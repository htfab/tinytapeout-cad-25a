VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_htfab_dg_dac
  CLASS BLOCK ;
  FOREIGN tt_um_htfab_dg_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.656000 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.150000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.227500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 32.000 5.000 34.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.000 5.000 100.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 65.000 5.000 67.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 35.000 5.000 37.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.000 5.000 103.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.000 5.000 70.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 38.000 5.000 40.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.000 5.000 106.000 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.000 5.000 73.000 220.760 ;
    END
  END VAPWR
  OBS
      LAYER nwell ;
        RECT 17.850 204.450 31.330 207.880 ;
        RECT 39.930 204.450 53.410 207.880 ;
        RECT 62.010 204.450 75.490 207.880 ;
        RECT 106.385 204.450 119.865 207.880 ;
      LAYER pwell ;
        RECT 17.850 204.200 18.780 204.205 ;
        RECT 39.930 204.200 40.860 204.205 ;
        RECT 62.010 204.200 62.940 204.205 ;
        RECT 106.385 204.200 107.315 204.205 ;
        RECT 17.850 201.420 31.330 204.200 ;
        RECT 39.930 201.420 53.410 204.200 ;
        RECT 62.010 201.420 75.490 204.200 ;
        RECT 106.385 201.420 119.865 204.200 ;
      LAYER nwell ;
        RECT 106.385 197.740 119.865 201.170 ;
      LAYER pwell ;
        RECT 106.385 197.490 107.315 197.495 ;
        RECT 106.385 194.710 119.865 197.490 ;
      LAYER nwell ;
        RECT 106.385 191.030 119.865 194.460 ;
      LAYER pwell ;
        RECT 106.385 190.780 107.315 190.785 ;
        RECT 106.385 188.000 119.865 190.780 ;
      LAYER nwell ;
        RECT 26.745 163.545 111.885 165.125 ;
        RECT 26.745 62.260 28.325 163.545 ;
      LAYER pwell ;
        RECT 42.530 160.765 96.450 163.545 ;
        RECT 55.080 160.760 56.010 160.765 ;
        RECT 68.560 160.760 69.490 160.765 ;
        RECT 82.040 160.760 82.970 160.765 ;
        RECT 95.520 160.760 96.450 160.765 ;
      LAYER nwell ;
        RECT 42.530 157.085 96.450 160.515 ;
      LAYER pwell ;
        RECT 35.965 154.135 38.750 155.065 ;
        RECT 35.965 140.085 38.745 154.135 ;
      LAYER nwell ;
        RECT 38.995 140.085 42.425 155.065 ;
      LAYER pwell ;
        RECT 42.675 154.135 45.460 155.065 ;
        RECT 42.675 140.085 45.455 154.135 ;
      LAYER nwell ;
        RECT 45.705 140.085 49.135 155.065 ;
      LAYER pwell ;
        RECT 49.385 154.135 52.170 155.065 ;
        RECT 49.385 140.085 52.165 154.135 ;
      LAYER nwell ;
        RECT 52.415 140.085 55.845 155.065 ;
      LAYER pwell ;
        RECT 56.095 154.135 58.880 155.065 ;
        RECT 56.095 140.085 58.875 154.135 ;
      LAYER nwell ;
        RECT 59.125 140.085 62.555 155.065 ;
      LAYER pwell ;
        RECT 62.805 154.135 65.590 155.065 ;
        RECT 62.805 140.085 65.585 154.135 ;
      LAYER nwell ;
        RECT 65.835 140.085 69.265 155.065 ;
      LAYER pwell ;
        RECT 69.515 154.135 72.300 155.065 ;
        RECT 69.515 140.085 72.295 154.135 ;
      LAYER nwell ;
        RECT 72.545 140.085 75.975 155.065 ;
      LAYER pwell ;
        RECT 76.225 154.135 79.010 155.065 ;
        RECT 76.225 140.085 79.005 154.135 ;
      LAYER nwell ;
        RECT 79.255 140.085 82.685 155.065 ;
      LAYER pwell ;
        RECT 82.935 154.135 85.720 155.065 ;
        RECT 82.935 140.085 85.715 154.135 ;
      LAYER nwell ;
        RECT 85.965 140.085 89.395 155.065 ;
      LAYER pwell ;
        RECT 89.645 154.135 92.430 155.065 ;
        RECT 89.645 140.085 92.425 154.135 ;
      LAYER nwell ;
        RECT 92.675 140.085 96.105 155.065 ;
      LAYER pwell ;
        RECT 96.355 154.135 99.140 155.065 ;
        RECT 96.355 140.085 99.135 154.135 ;
      LAYER nwell ;
        RECT 99.385 140.085 102.815 155.065 ;
      LAYER pwell ;
        RECT 55.505 128.635 83.155 133.155 ;
      LAYER nwell ;
        RECT 55.505 122.775 83.205 128.385 ;
      LAYER pwell ;
        RECT 54.800 107.110 83.910 122.220 ;
      LAYER nwell ;
        RECT 55.505 100.945 83.205 106.555 ;
      LAYER pwell ;
        RECT 55.555 96.175 83.205 100.695 ;
      LAYER nwell ;
        RECT 30.325 88.645 108.305 92.075 ;
      LAYER pwell ;
        RECT 30.325 88.395 31.255 88.400 ;
        RECT 30.325 85.615 108.305 88.395 ;
      LAYER nwell ;
        RECT 35.990 64.260 39.420 79.240 ;
      LAYER pwell ;
        RECT 39.670 65.190 42.450 79.240 ;
        RECT 39.665 64.260 42.450 65.190 ;
      LAYER nwell ;
        RECT 42.700 64.260 46.130 79.240 ;
      LAYER pwell ;
        RECT 46.380 65.190 49.160 79.240 ;
        RECT 46.375 64.260 49.160 65.190 ;
      LAYER nwell ;
        RECT 49.410 64.260 52.840 79.240 ;
      LAYER pwell ;
        RECT 53.090 65.190 55.870 79.240 ;
        RECT 53.085 64.260 55.870 65.190 ;
      LAYER nwell ;
        RECT 56.120 64.260 59.550 79.240 ;
      LAYER pwell ;
        RECT 59.800 65.190 62.580 79.240 ;
        RECT 59.795 64.260 62.580 65.190 ;
      LAYER nwell ;
        RECT 62.830 64.260 66.260 79.240 ;
      LAYER pwell ;
        RECT 66.510 65.190 69.290 79.240 ;
        RECT 66.505 64.260 69.290 65.190 ;
      LAYER nwell ;
        RECT 69.540 64.260 72.970 79.240 ;
      LAYER pwell ;
        RECT 73.220 65.190 76.000 79.240 ;
        RECT 73.215 64.260 76.000 65.190 ;
      LAYER nwell ;
        RECT 76.250 64.260 79.680 79.240 ;
      LAYER pwell ;
        RECT 79.930 65.190 82.710 79.240 ;
        RECT 79.925 64.260 82.710 65.190 ;
      LAYER nwell ;
        RECT 82.960 64.260 86.390 79.240 ;
      LAYER pwell ;
        RECT 86.640 65.190 89.420 79.240 ;
        RECT 86.635 64.260 89.420 65.190 ;
      LAYER nwell ;
        RECT 89.670 64.260 93.100 79.240 ;
      LAYER pwell ;
        RECT 93.350 65.190 96.130 79.240 ;
        RECT 93.345 64.260 96.130 65.190 ;
      LAYER nwell ;
        RECT 96.380 64.260 99.810 79.240 ;
      LAYER pwell ;
        RECT 100.060 65.190 102.840 79.240 ;
        RECT 100.055 64.260 102.840 65.190 ;
      LAYER nwell ;
        RECT 110.305 62.260 111.885 163.545 ;
        RECT 26.745 60.680 111.885 62.260 ;
      LAYER li1 ;
        RECT 18.240 207.320 30.940 207.490 ;
        RECT 18.240 205.100 18.410 207.320 ;
        RECT 19.090 206.900 19.590 207.070 ;
        RECT 20.590 206.900 21.090 207.070 ;
        RECT 22.090 206.900 22.590 207.070 ;
        RECT 23.590 206.900 24.090 207.070 ;
        RECT 25.090 206.900 25.590 207.070 ;
        RECT 26.590 206.900 27.090 207.070 ;
        RECT 28.090 206.900 28.590 207.070 ;
        RECT 29.590 206.900 30.090 207.070 ;
        RECT 18.800 205.645 18.970 206.685 ;
        RECT 19.710 205.645 19.880 206.685 ;
        RECT 20.300 205.645 20.470 206.685 ;
        RECT 21.210 205.645 21.380 206.685 ;
        RECT 21.800 205.645 21.970 206.685 ;
        RECT 22.710 205.645 22.880 206.685 ;
        RECT 23.300 205.645 23.470 206.685 ;
        RECT 24.210 205.645 24.380 206.685 ;
        RECT 24.800 205.645 24.970 206.685 ;
        RECT 25.710 205.645 25.880 206.685 ;
        RECT 26.300 205.645 26.470 206.685 ;
        RECT 27.210 205.645 27.380 206.685 ;
        RECT 27.800 205.645 27.970 206.685 ;
        RECT 28.710 205.645 28.880 206.685 ;
        RECT 29.300 205.645 29.470 206.685 ;
        RECT 30.210 205.645 30.380 206.685 ;
        RECT 19.090 205.260 19.590 205.430 ;
        RECT 20.590 205.260 21.090 205.430 ;
        RECT 22.090 205.260 22.590 205.430 ;
        RECT 23.590 205.260 24.090 205.430 ;
        RECT 25.090 205.260 25.590 205.430 ;
        RECT 26.590 205.260 27.090 205.430 ;
        RECT 28.090 205.260 28.590 205.430 ;
        RECT 29.590 205.260 30.090 205.430 ;
        RECT 30.770 205.100 30.940 207.320 ;
        RECT 40.320 207.320 53.020 207.490 ;
        RECT 40.320 205.100 40.490 207.320 ;
        RECT 41.170 206.900 41.670 207.070 ;
        RECT 42.670 206.900 43.170 207.070 ;
        RECT 44.170 206.900 44.670 207.070 ;
        RECT 45.670 206.900 46.170 207.070 ;
        RECT 47.170 206.900 47.670 207.070 ;
        RECT 48.670 206.900 49.170 207.070 ;
        RECT 50.170 206.900 50.670 207.070 ;
        RECT 51.670 206.900 52.170 207.070 ;
        RECT 40.880 205.645 41.050 206.685 ;
        RECT 41.790 205.645 41.960 206.685 ;
        RECT 42.380 205.645 42.550 206.685 ;
        RECT 43.290 205.645 43.460 206.685 ;
        RECT 43.880 205.645 44.050 206.685 ;
        RECT 44.790 205.645 44.960 206.685 ;
        RECT 45.380 205.645 45.550 206.685 ;
        RECT 46.290 205.645 46.460 206.685 ;
        RECT 46.880 205.645 47.050 206.685 ;
        RECT 47.790 205.645 47.960 206.685 ;
        RECT 48.380 205.645 48.550 206.685 ;
        RECT 49.290 205.645 49.460 206.685 ;
        RECT 49.880 205.645 50.050 206.685 ;
        RECT 50.790 205.645 50.960 206.685 ;
        RECT 51.380 205.645 51.550 206.685 ;
        RECT 52.290 205.645 52.460 206.685 ;
        RECT 41.170 205.260 41.670 205.430 ;
        RECT 42.670 205.260 43.170 205.430 ;
        RECT 44.170 205.260 44.670 205.430 ;
        RECT 45.670 205.260 46.170 205.430 ;
        RECT 47.170 205.260 47.670 205.430 ;
        RECT 48.670 205.260 49.170 205.430 ;
        RECT 50.170 205.260 50.670 205.430 ;
        RECT 51.670 205.260 52.170 205.430 ;
        RECT 52.850 205.100 53.020 207.320 ;
        RECT 62.400 207.320 75.100 207.490 ;
        RECT 62.400 205.100 62.570 207.320 ;
        RECT 63.250 206.900 63.750 207.070 ;
        RECT 64.750 206.900 65.250 207.070 ;
        RECT 66.250 206.900 66.750 207.070 ;
        RECT 67.750 206.900 68.250 207.070 ;
        RECT 69.250 206.900 69.750 207.070 ;
        RECT 70.750 206.900 71.250 207.070 ;
        RECT 72.250 206.900 72.750 207.070 ;
        RECT 73.750 206.900 74.250 207.070 ;
        RECT 62.960 205.645 63.130 206.685 ;
        RECT 63.870 205.645 64.040 206.685 ;
        RECT 64.460 205.645 64.630 206.685 ;
        RECT 65.370 205.645 65.540 206.685 ;
        RECT 65.960 205.645 66.130 206.685 ;
        RECT 66.870 205.645 67.040 206.685 ;
        RECT 67.460 205.645 67.630 206.685 ;
        RECT 68.370 205.645 68.540 206.685 ;
        RECT 68.960 205.645 69.130 206.685 ;
        RECT 69.870 205.645 70.040 206.685 ;
        RECT 70.460 205.645 70.630 206.685 ;
        RECT 71.370 205.645 71.540 206.685 ;
        RECT 71.960 205.645 72.130 206.685 ;
        RECT 72.870 205.645 73.040 206.685 ;
        RECT 73.460 205.645 73.630 206.685 ;
        RECT 74.370 205.645 74.540 206.685 ;
        RECT 63.250 205.260 63.750 205.430 ;
        RECT 64.750 205.260 65.250 205.430 ;
        RECT 66.250 205.260 66.750 205.430 ;
        RECT 67.750 205.260 68.250 205.430 ;
        RECT 69.250 205.260 69.750 205.430 ;
        RECT 70.750 205.260 71.250 205.430 ;
        RECT 72.250 205.260 72.750 205.430 ;
        RECT 73.750 205.260 74.250 205.430 ;
        RECT 74.930 205.100 75.100 207.320 ;
        RECT 106.775 207.320 119.475 207.490 ;
        RECT 106.775 205.100 106.945 207.320 ;
        RECT 107.625 206.900 108.125 207.070 ;
        RECT 109.125 206.900 109.625 207.070 ;
        RECT 110.625 206.900 111.125 207.070 ;
        RECT 112.125 206.900 112.625 207.070 ;
        RECT 113.625 206.900 114.125 207.070 ;
        RECT 115.125 206.900 115.625 207.070 ;
        RECT 116.625 206.900 117.125 207.070 ;
        RECT 118.125 206.900 118.625 207.070 ;
        RECT 107.335 205.645 107.505 206.685 ;
        RECT 108.245 205.645 108.415 206.685 ;
        RECT 108.835 205.645 109.005 206.685 ;
        RECT 109.745 205.645 109.915 206.685 ;
        RECT 110.335 205.645 110.505 206.685 ;
        RECT 111.245 205.645 111.415 206.685 ;
        RECT 111.835 205.645 112.005 206.685 ;
        RECT 112.745 205.645 112.915 206.685 ;
        RECT 113.335 205.645 113.505 206.685 ;
        RECT 114.245 205.645 114.415 206.685 ;
        RECT 114.835 205.645 115.005 206.685 ;
        RECT 115.745 205.645 115.915 206.685 ;
        RECT 116.335 205.645 116.505 206.685 ;
        RECT 117.245 205.645 117.415 206.685 ;
        RECT 117.835 205.645 118.005 206.685 ;
        RECT 118.745 205.645 118.915 206.685 ;
        RECT 107.625 205.260 108.125 205.430 ;
        RECT 109.125 205.260 109.625 205.430 ;
        RECT 110.625 205.260 111.125 205.430 ;
        RECT 112.125 205.260 112.625 205.430 ;
        RECT 113.625 205.260 114.125 205.430 ;
        RECT 115.125 205.260 115.625 205.430 ;
        RECT 116.625 205.260 117.125 205.430 ;
        RECT 118.125 205.260 118.625 205.430 ;
        RECT 18.240 205.010 18.850 205.100 ;
        RECT 30.770 205.010 31.330 205.100 ;
        RECT 18.240 204.840 31.330 205.010 ;
        RECT 40.320 205.010 40.930 205.100 ;
        RECT 52.850 205.010 53.410 205.100 ;
        RECT 40.320 204.840 53.410 205.010 ;
        RECT 62.400 205.010 63.010 205.100 ;
        RECT 74.930 205.010 75.490 205.100 ;
        RECT 62.400 204.840 75.490 205.010 ;
        RECT 18.350 204.750 18.850 204.840 ;
        RECT 30.770 204.750 31.330 204.840 ;
        RECT 40.430 204.750 40.930 204.840 ;
        RECT 52.850 204.750 53.410 204.840 ;
        RECT 62.510 204.750 63.010 204.840 ;
        RECT 74.930 204.750 75.490 204.840 ;
        RECT 106.370 205.010 106.945 205.100 ;
        RECT 119.305 205.100 119.475 207.320 ;
        RECT 119.305 205.010 119.945 205.100 ;
        RECT 106.370 204.840 119.945 205.010 ;
        RECT 106.370 204.750 106.870 204.840 ;
        RECT 119.445 204.750 119.945 204.840 ;
        RECT 18.140 203.960 18.850 204.050 ;
        RECT 30.830 203.960 31.330 204.050 ;
        RECT 18.140 203.790 31.330 203.960 ;
        RECT 18.140 203.700 18.850 203.790 ;
        RECT 30.830 203.700 31.330 203.790 ;
        RECT 40.220 203.960 40.930 204.050 ;
        RECT 52.910 203.960 53.410 204.050 ;
        RECT 40.220 203.790 53.410 203.960 ;
        RECT 40.220 203.700 40.930 203.790 ;
        RECT 52.910 203.700 53.410 203.790 ;
        RECT 62.300 203.960 63.010 204.050 ;
        RECT 74.990 203.960 75.490 204.050 ;
        RECT 62.300 203.790 75.490 203.960 ;
        RECT 62.300 203.700 63.010 203.790 ;
        RECT 74.990 203.700 75.490 203.790 ;
        RECT 106.370 203.960 106.870 204.050 ;
        RECT 119.445 203.960 119.945 204.050 ;
        RECT 106.370 203.790 119.945 203.960 ;
        RECT 106.370 203.700 106.870 203.790 ;
        RECT 119.445 203.700 119.945 203.790 ;
        RECT 18.140 201.830 18.310 203.700 ;
        RECT 19.090 203.325 19.590 203.495 ;
        RECT 20.590 203.325 21.090 203.495 ;
        RECT 22.090 203.325 22.590 203.495 ;
        RECT 23.590 203.325 24.090 203.495 ;
        RECT 25.090 203.325 25.590 203.495 ;
        RECT 26.590 203.325 27.090 203.495 ;
        RECT 28.090 203.325 28.590 203.495 ;
        RECT 29.590 203.325 30.090 203.495 ;
        RECT 18.800 202.465 18.970 203.155 ;
        RECT 19.710 202.465 19.880 203.155 ;
        RECT 20.300 202.465 20.470 203.155 ;
        RECT 21.210 202.465 21.380 203.155 ;
        RECT 21.800 202.465 21.970 203.155 ;
        RECT 22.710 202.465 22.880 203.155 ;
        RECT 23.300 202.465 23.470 203.155 ;
        RECT 24.210 202.465 24.380 203.155 ;
        RECT 24.800 202.465 24.970 203.155 ;
        RECT 25.710 202.465 25.880 203.155 ;
        RECT 26.300 202.465 26.470 203.155 ;
        RECT 27.210 202.465 27.380 203.155 ;
        RECT 27.800 202.465 27.970 203.155 ;
        RECT 28.710 202.465 28.880 203.155 ;
        RECT 29.300 202.465 29.470 203.155 ;
        RECT 30.210 202.465 30.380 203.155 ;
        RECT 19.090 202.125 19.590 202.295 ;
        RECT 20.590 202.125 21.090 202.295 ;
        RECT 22.090 202.125 22.590 202.295 ;
        RECT 23.590 202.125 24.090 202.295 ;
        RECT 25.090 202.125 25.590 202.295 ;
        RECT 26.590 202.125 27.090 202.295 ;
        RECT 28.090 202.125 28.590 202.295 ;
        RECT 29.590 202.125 30.090 202.295 ;
        RECT 30.920 201.830 31.090 203.700 ;
        RECT 18.140 201.660 31.090 201.830 ;
        RECT 40.220 201.830 40.390 203.700 ;
        RECT 41.170 203.325 41.670 203.495 ;
        RECT 42.670 203.325 43.170 203.495 ;
        RECT 44.170 203.325 44.670 203.495 ;
        RECT 45.670 203.325 46.170 203.495 ;
        RECT 47.170 203.325 47.670 203.495 ;
        RECT 48.670 203.325 49.170 203.495 ;
        RECT 50.170 203.325 50.670 203.495 ;
        RECT 51.670 203.325 52.170 203.495 ;
        RECT 40.880 202.465 41.050 203.155 ;
        RECT 41.790 202.465 41.960 203.155 ;
        RECT 42.380 202.465 42.550 203.155 ;
        RECT 43.290 202.465 43.460 203.155 ;
        RECT 43.880 202.465 44.050 203.155 ;
        RECT 44.790 202.465 44.960 203.155 ;
        RECT 45.380 202.465 45.550 203.155 ;
        RECT 46.290 202.465 46.460 203.155 ;
        RECT 46.880 202.465 47.050 203.155 ;
        RECT 47.790 202.465 47.960 203.155 ;
        RECT 48.380 202.465 48.550 203.155 ;
        RECT 49.290 202.465 49.460 203.155 ;
        RECT 49.880 202.465 50.050 203.155 ;
        RECT 50.790 202.465 50.960 203.155 ;
        RECT 51.380 202.465 51.550 203.155 ;
        RECT 52.290 202.465 52.460 203.155 ;
        RECT 41.170 202.125 41.670 202.295 ;
        RECT 42.670 202.125 43.170 202.295 ;
        RECT 44.170 202.125 44.670 202.295 ;
        RECT 45.670 202.125 46.170 202.295 ;
        RECT 47.170 202.125 47.670 202.295 ;
        RECT 48.670 202.125 49.170 202.295 ;
        RECT 50.170 202.125 50.670 202.295 ;
        RECT 51.670 202.125 52.170 202.295 ;
        RECT 53.000 201.830 53.170 203.700 ;
        RECT 40.220 201.660 53.170 201.830 ;
        RECT 62.300 201.830 62.470 203.700 ;
        RECT 63.250 203.325 63.750 203.495 ;
        RECT 64.750 203.325 65.250 203.495 ;
        RECT 66.250 203.325 66.750 203.495 ;
        RECT 67.750 203.325 68.250 203.495 ;
        RECT 69.250 203.325 69.750 203.495 ;
        RECT 70.750 203.325 71.250 203.495 ;
        RECT 72.250 203.325 72.750 203.495 ;
        RECT 73.750 203.325 74.250 203.495 ;
        RECT 62.960 202.465 63.130 203.155 ;
        RECT 63.870 202.465 64.040 203.155 ;
        RECT 64.460 202.465 64.630 203.155 ;
        RECT 65.370 202.465 65.540 203.155 ;
        RECT 65.960 202.465 66.130 203.155 ;
        RECT 66.870 202.465 67.040 203.155 ;
        RECT 67.460 202.465 67.630 203.155 ;
        RECT 68.370 202.465 68.540 203.155 ;
        RECT 68.960 202.465 69.130 203.155 ;
        RECT 69.870 202.465 70.040 203.155 ;
        RECT 70.460 202.465 70.630 203.155 ;
        RECT 71.370 202.465 71.540 203.155 ;
        RECT 71.960 202.465 72.130 203.155 ;
        RECT 72.870 202.465 73.040 203.155 ;
        RECT 73.460 202.465 73.630 203.155 ;
        RECT 74.370 202.465 74.540 203.155 ;
        RECT 63.250 202.125 63.750 202.295 ;
        RECT 64.750 202.125 65.250 202.295 ;
        RECT 66.250 202.125 66.750 202.295 ;
        RECT 67.750 202.125 68.250 202.295 ;
        RECT 69.250 202.125 69.750 202.295 ;
        RECT 70.750 202.125 71.250 202.295 ;
        RECT 72.250 202.125 72.750 202.295 ;
        RECT 73.750 202.125 74.250 202.295 ;
        RECT 75.080 201.830 75.250 203.700 ;
        RECT 62.300 201.660 75.250 201.830 ;
        RECT 106.675 201.830 106.845 203.700 ;
        RECT 107.625 203.325 108.125 203.495 ;
        RECT 109.125 203.325 109.625 203.495 ;
        RECT 110.625 203.325 111.125 203.495 ;
        RECT 112.125 203.325 112.625 203.495 ;
        RECT 113.625 203.325 114.125 203.495 ;
        RECT 115.125 203.325 115.625 203.495 ;
        RECT 116.625 203.325 117.125 203.495 ;
        RECT 118.125 203.325 118.625 203.495 ;
        RECT 107.335 202.465 107.505 203.155 ;
        RECT 108.245 202.465 108.415 203.155 ;
        RECT 108.835 202.465 109.005 203.155 ;
        RECT 109.745 202.465 109.915 203.155 ;
        RECT 110.335 202.465 110.505 203.155 ;
        RECT 111.245 202.465 111.415 203.155 ;
        RECT 111.835 202.465 112.005 203.155 ;
        RECT 112.745 202.465 112.915 203.155 ;
        RECT 113.335 202.465 113.505 203.155 ;
        RECT 114.245 202.465 114.415 203.155 ;
        RECT 114.835 202.465 115.005 203.155 ;
        RECT 115.745 202.465 115.915 203.155 ;
        RECT 116.335 202.465 116.505 203.155 ;
        RECT 117.245 202.465 117.415 203.155 ;
        RECT 117.835 202.465 118.005 203.155 ;
        RECT 118.745 202.465 118.915 203.155 ;
        RECT 107.625 202.125 108.125 202.295 ;
        RECT 109.125 202.125 109.625 202.295 ;
        RECT 110.625 202.125 111.125 202.295 ;
        RECT 112.125 202.125 112.625 202.295 ;
        RECT 113.625 202.125 114.125 202.295 ;
        RECT 115.125 202.125 115.625 202.295 ;
        RECT 116.625 202.125 117.125 202.295 ;
        RECT 118.125 202.125 118.625 202.295 ;
        RECT 119.455 201.830 119.625 203.700 ;
        RECT 106.675 201.660 119.625 201.830 ;
        RECT 106.775 200.610 119.475 200.780 ;
        RECT 106.775 198.390 106.945 200.610 ;
        RECT 107.625 200.190 108.125 200.360 ;
        RECT 109.125 200.190 109.625 200.360 ;
        RECT 110.625 200.190 111.125 200.360 ;
        RECT 112.125 200.190 112.625 200.360 ;
        RECT 113.625 200.190 114.125 200.360 ;
        RECT 115.125 200.190 115.625 200.360 ;
        RECT 116.625 200.190 117.125 200.360 ;
        RECT 118.125 200.190 118.625 200.360 ;
        RECT 107.335 198.935 107.505 199.975 ;
        RECT 108.245 198.935 108.415 199.975 ;
        RECT 108.835 198.935 109.005 199.975 ;
        RECT 109.745 198.935 109.915 199.975 ;
        RECT 110.335 198.935 110.505 199.975 ;
        RECT 111.245 198.935 111.415 199.975 ;
        RECT 111.835 198.935 112.005 199.975 ;
        RECT 112.745 198.935 112.915 199.975 ;
        RECT 113.335 198.935 113.505 199.975 ;
        RECT 114.245 198.935 114.415 199.975 ;
        RECT 114.835 198.935 115.005 199.975 ;
        RECT 115.745 198.935 115.915 199.975 ;
        RECT 116.335 198.935 116.505 199.975 ;
        RECT 117.245 198.935 117.415 199.975 ;
        RECT 117.835 198.935 118.005 199.975 ;
        RECT 118.745 198.935 118.915 199.975 ;
        RECT 107.625 198.550 108.125 198.720 ;
        RECT 109.125 198.550 109.625 198.720 ;
        RECT 110.625 198.550 111.125 198.720 ;
        RECT 112.125 198.550 112.625 198.720 ;
        RECT 113.625 198.550 114.125 198.720 ;
        RECT 115.125 198.550 115.625 198.720 ;
        RECT 116.625 198.550 117.125 198.720 ;
        RECT 118.125 198.550 118.625 198.720 ;
        RECT 106.370 198.300 106.945 198.390 ;
        RECT 119.305 198.390 119.475 200.610 ;
        RECT 119.305 198.300 119.945 198.390 ;
        RECT 106.370 198.130 119.945 198.300 ;
        RECT 106.370 198.040 106.870 198.130 ;
        RECT 119.445 198.040 119.945 198.130 ;
        RECT 106.370 197.250 106.870 197.340 ;
        RECT 119.445 197.250 119.945 197.340 ;
        RECT 106.370 197.080 119.945 197.250 ;
        RECT 106.370 196.990 106.870 197.080 ;
        RECT 119.445 196.990 119.945 197.080 ;
        RECT 106.675 195.120 106.845 196.990 ;
        RECT 107.625 196.615 108.125 196.785 ;
        RECT 109.125 196.615 109.625 196.785 ;
        RECT 110.625 196.615 111.125 196.785 ;
        RECT 112.125 196.615 112.625 196.785 ;
        RECT 113.625 196.615 114.125 196.785 ;
        RECT 115.125 196.615 115.625 196.785 ;
        RECT 116.625 196.615 117.125 196.785 ;
        RECT 118.125 196.615 118.625 196.785 ;
        RECT 107.335 195.755 107.505 196.445 ;
        RECT 108.245 195.755 108.415 196.445 ;
        RECT 108.835 195.755 109.005 196.445 ;
        RECT 109.745 195.755 109.915 196.445 ;
        RECT 110.335 195.755 110.505 196.445 ;
        RECT 111.245 195.755 111.415 196.445 ;
        RECT 111.835 195.755 112.005 196.445 ;
        RECT 112.745 195.755 112.915 196.445 ;
        RECT 113.335 195.755 113.505 196.445 ;
        RECT 114.245 195.755 114.415 196.445 ;
        RECT 114.835 195.755 115.005 196.445 ;
        RECT 115.745 195.755 115.915 196.445 ;
        RECT 116.335 195.755 116.505 196.445 ;
        RECT 117.245 195.755 117.415 196.445 ;
        RECT 117.835 195.755 118.005 196.445 ;
        RECT 118.745 195.755 118.915 196.445 ;
        RECT 107.625 195.415 108.125 195.585 ;
        RECT 109.125 195.415 109.625 195.585 ;
        RECT 110.625 195.415 111.125 195.585 ;
        RECT 112.125 195.415 112.625 195.585 ;
        RECT 113.625 195.415 114.125 195.585 ;
        RECT 115.125 195.415 115.625 195.585 ;
        RECT 116.625 195.415 117.125 195.585 ;
        RECT 118.125 195.415 118.625 195.585 ;
        RECT 119.455 195.120 119.625 196.990 ;
        RECT 106.675 194.950 119.625 195.120 ;
        RECT 106.775 193.900 119.475 194.070 ;
        RECT 106.775 191.680 106.945 193.900 ;
        RECT 107.625 193.480 108.125 193.650 ;
        RECT 109.125 193.480 109.625 193.650 ;
        RECT 110.625 193.480 111.125 193.650 ;
        RECT 112.125 193.480 112.625 193.650 ;
        RECT 113.625 193.480 114.125 193.650 ;
        RECT 115.125 193.480 115.625 193.650 ;
        RECT 116.625 193.480 117.125 193.650 ;
        RECT 118.125 193.480 118.625 193.650 ;
        RECT 107.335 192.225 107.505 193.265 ;
        RECT 108.245 192.225 108.415 193.265 ;
        RECT 108.835 192.225 109.005 193.265 ;
        RECT 109.745 192.225 109.915 193.265 ;
        RECT 110.335 192.225 110.505 193.265 ;
        RECT 111.245 192.225 111.415 193.265 ;
        RECT 111.835 192.225 112.005 193.265 ;
        RECT 112.745 192.225 112.915 193.265 ;
        RECT 113.335 192.225 113.505 193.265 ;
        RECT 114.245 192.225 114.415 193.265 ;
        RECT 114.835 192.225 115.005 193.265 ;
        RECT 115.745 192.225 115.915 193.265 ;
        RECT 116.335 192.225 116.505 193.265 ;
        RECT 117.245 192.225 117.415 193.265 ;
        RECT 117.835 192.225 118.005 193.265 ;
        RECT 118.745 192.225 118.915 193.265 ;
        RECT 107.625 191.840 108.125 192.010 ;
        RECT 109.125 191.840 109.625 192.010 ;
        RECT 110.625 191.840 111.125 192.010 ;
        RECT 112.125 191.840 112.625 192.010 ;
        RECT 113.625 191.840 114.125 192.010 ;
        RECT 115.125 191.840 115.625 192.010 ;
        RECT 116.625 191.840 117.125 192.010 ;
        RECT 118.125 191.840 118.625 192.010 ;
        RECT 106.370 191.590 106.945 191.680 ;
        RECT 119.305 191.680 119.475 193.900 ;
        RECT 119.305 191.590 119.945 191.680 ;
        RECT 106.370 191.420 119.945 191.590 ;
        RECT 106.370 191.330 106.870 191.420 ;
        RECT 119.445 191.330 119.945 191.420 ;
        RECT 106.370 190.540 106.870 190.630 ;
        RECT 119.445 190.540 119.945 190.630 ;
        RECT 106.370 190.370 119.945 190.540 ;
        RECT 106.370 190.280 106.870 190.370 ;
        RECT 119.445 190.280 119.945 190.370 ;
        RECT 106.675 188.410 106.845 190.280 ;
        RECT 107.625 189.905 108.125 190.075 ;
        RECT 109.125 189.905 109.625 190.075 ;
        RECT 110.625 189.905 111.125 190.075 ;
        RECT 112.125 189.905 112.625 190.075 ;
        RECT 113.625 189.905 114.125 190.075 ;
        RECT 115.125 189.905 115.625 190.075 ;
        RECT 116.625 189.905 117.125 190.075 ;
        RECT 118.125 189.905 118.625 190.075 ;
        RECT 107.335 189.045 107.505 189.735 ;
        RECT 108.245 189.045 108.415 189.735 ;
        RECT 108.835 189.045 109.005 189.735 ;
        RECT 109.745 189.045 109.915 189.735 ;
        RECT 110.335 189.045 110.505 189.735 ;
        RECT 111.245 189.045 111.415 189.735 ;
        RECT 111.835 189.045 112.005 189.735 ;
        RECT 112.745 189.045 112.915 189.735 ;
        RECT 113.335 189.045 113.505 189.735 ;
        RECT 114.245 189.045 114.415 189.735 ;
        RECT 114.835 189.045 115.005 189.735 ;
        RECT 115.745 189.045 115.915 189.735 ;
        RECT 116.335 189.045 116.505 189.735 ;
        RECT 117.245 189.045 117.415 189.735 ;
        RECT 117.835 189.045 118.005 189.735 ;
        RECT 118.745 189.045 118.915 189.735 ;
        RECT 107.625 188.705 108.125 188.875 ;
        RECT 109.125 188.705 109.625 188.875 ;
        RECT 110.625 188.705 111.125 188.875 ;
        RECT 112.125 188.705 112.625 188.875 ;
        RECT 113.625 188.705 114.125 188.875 ;
        RECT 115.125 188.705 115.625 188.875 ;
        RECT 116.625 188.705 117.125 188.875 ;
        RECT 118.125 188.705 118.625 188.875 ;
        RECT 119.455 188.410 119.625 190.280 ;
        RECT 106.675 188.240 119.625 188.410 ;
        RECT 27.180 164.520 111.450 164.690 ;
        RECT 27.180 61.285 27.350 164.520 ;
        RECT 42.770 163.135 55.720 163.305 ;
        RECT 42.770 161.175 42.940 163.135 ;
        RECT 43.770 162.670 44.270 162.840 ;
        RECT 45.270 162.670 45.770 162.840 ;
        RECT 46.770 162.670 47.270 162.840 ;
        RECT 48.270 162.670 48.770 162.840 ;
        RECT 49.770 162.670 50.270 162.840 ;
        RECT 51.270 162.670 51.770 162.840 ;
        RECT 52.770 162.670 53.270 162.840 ;
        RECT 54.270 162.670 54.770 162.840 ;
        RECT 43.480 161.810 43.650 162.500 ;
        RECT 44.390 161.810 44.560 162.500 ;
        RECT 44.980 161.810 45.150 162.500 ;
        RECT 45.890 161.810 46.060 162.500 ;
        RECT 46.480 161.810 46.650 162.500 ;
        RECT 47.390 161.810 47.560 162.500 ;
        RECT 47.980 161.810 48.150 162.500 ;
        RECT 48.890 161.810 49.060 162.500 ;
        RECT 49.480 161.810 49.650 162.500 ;
        RECT 50.390 161.810 50.560 162.500 ;
        RECT 50.980 161.810 51.150 162.500 ;
        RECT 51.890 161.810 52.060 162.500 ;
        RECT 52.480 161.810 52.650 162.500 ;
        RECT 53.390 161.810 53.560 162.500 ;
        RECT 53.980 161.810 54.150 162.500 ;
        RECT 54.890 161.810 55.060 162.500 ;
        RECT 43.770 161.470 44.270 161.640 ;
        RECT 45.270 161.470 45.770 161.640 ;
        RECT 46.770 161.470 47.270 161.640 ;
        RECT 48.270 161.470 48.770 161.640 ;
        RECT 49.770 161.470 50.270 161.640 ;
        RECT 51.270 161.470 51.770 161.640 ;
        RECT 52.770 161.470 53.270 161.640 ;
        RECT 54.270 161.470 54.770 161.640 ;
        RECT 55.550 161.175 55.720 163.135 ;
        RECT 42.770 161.005 55.720 161.175 ;
        RECT 56.250 163.135 69.200 163.305 ;
        RECT 56.250 161.175 56.420 163.135 ;
        RECT 57.250 162.670 57.750 162.840 ;
        RECT 58.750 162.670 59.250 162.840 ;
        RECT 60.250 162.670 60.750 162.840 ;
        RECT 61.750 162.670 62.250 162.840 ;
        RECT 63.250 162.670 63.750 162.840 ;
        RECT 64.750 162.670 65.250 162.840 ;
        RECT 66.250 162.670 66.750 162.840 ;
        RECT 67.750 162.670 68.250 162.840 ;
        RECT 56.960 161.810 57.130 162.500 ;
        RECT 57.870 161.810 58.040 162.500 ;
        RECT 58.460 161.810 58.630 162.500 ;
        RECT 59.370 161.810 59.540 162.500 ;
        RECT 59.960 161.810 60.130 162.500 ;
        RECT 60.870 161.810 61.040 162.500 ;
        RECT 61.460 161.810 61.630 162.500 ;
        RECT 62.370 161.810 62.540 162.500 ;
        RECT 62.960 161.810 63.130 162.500 ;
        RECT 63.870 161.810 64.040 162.500 ;
        RECT 64.460 161.810 64.630 162.500 ;
        RECT 65.370 161.810 65.540 162.500 ;
        RECT 65.960 161.810 66.130 162.500 ;
        RECT 66.870 161.810 67.040 162.500 ;
        RECT 67.460 161.810 67.630 162.500 ;
        RECT 68.370 161.810 68.540 162.500 ;
        RECT 57.250 161.470 57.750 161.640 ;
        RECT 58.750 161.470 59.250 161.640 ;
        RECT 60.250 161.470 60.750 161.640 ;
        RECT 61.750 161.470 62.250 161.640 ;
        RECT 63.250 161.470 63.750 161.640 ;
        RECT 64.750 161.470 65.250 161.640 ;
        RECT 66.250 161.470 66.750 161.640 ;
        RECT 67.750 161.470 68.250 161.640 ;
        RECT 69.030 161.175 69.200 163.135 ;
        RECT 56.250 161.005 69.200 161.175 ;
        RECT 69.730 163.135 82.680 163.305 ;
        RECT 69.730 161.175 69.900 163.135 ;
        RECT 70.730 162.670 71.230 162.840 ;
        RECT 72.230 162.670 72.730 162.840 ;
        RECT 73.730 162.670 74.230 162.840 ;
        RECT 75.230 162.670 75.730 162.840 ;
        RECT 76.730 162.670 77.230 162.840 ;
        RECT 78.230 162.670 78.730 162.840 ;
        RECT 79.730 162.670 80.230 162.840 ;
        RECT 81.230 162.670 81.730 162.840 ;
        RECT 70.440 161.810 70.610 162.500 ;
        RECT 71.350 161.810 71.520 162.500 ;
        RECT 71.940 161.810 72.110 162.500 ;
        RECT 72.850 161.810 73.020 162.500 ;
        RECT 73.440 161.810 73.610 162.500 ;
        RECT 74.350 161.810 74.520 162.500 ;
        RECT 74.940 161.810 75.110 162.500 ;
        RECT 75.850 161.810 76.020 162.500 ;
        RECT 76.440 161.810 76.610 162.500 ;
        RECT 77.350 161.810 77.520 162.500 ;
        RECT 77.940 161.810 78.110 162.500 ;
        RECT 78.850 161.810 79.020 162.500 ;
        RECT 79.440 161.810 79.610 162.500 ;
        RECT 80.350 161.810 80.520 162.500 ;
        RECT 80.940 161.810 81.110 162.500 ;
        RECT 81.850 161.810 82.020 162.500 ;
        RECT 70.730 161.470 71.230 161.640 ;
        RECT 72.230 161.470 72.730 161.640 ;
        RECT 73.730 161.470 74.230 161.640 ;
        RECT 75.230 161.470 75.730 161.640 ;
        RECT 76.730 161.470 77.230 161.640 ;
        RECT 78.230 161.470 78.730 161.640 ;
        RECT 79.730 161.470 80.230 161.640 ;
        RECT 81.230 161.470 81.730 161.640 ;
        RECT 82.510 161.175 82.680 163.135 ;
        RECT 69.730 161.005 82.680 161.175 ;
        RECT 83.210 163.135 96.160 163.305 ;
        RECT 83.210 161.175 83.380 163.135 ;
        RECT 84.210 162.670 84.710 162.840 ;
        RECT 85.710 162.670 86.210 162.840 ;
        RECT 87.210 162.670 87.710 162.840 ;
        RECT 88.710 162.670 89.210 162.840 ;
        RECT 90.210 162.670 90.710 162.840 ;
        RECT 91.710 162.670 92.210 162.840 ;
        RECT 93.210 162.670 93.710 162.840 ;
        RECT 94.710 162.670 95.210 162.840 ;
        RECT 83.920 161.810 84.090 162.500 ;
        RECT 84.830 161.810 85.000 162.500 ;
        RECT 85.420 161.810 85.590 162.500 ;
        RECT 86.330 161.810 86.500 162.500 ;
        RECT 86.920 161.810 87.090 162.500 ;
        RECT 87.830 161.810 88.000 162.500 ;
        RECT 88.420 161.810 88.590 162.500 ;
        RECT 89.330 161.810 89.500 162.500 ;
        RECT 89.920 161.810 90.090 162.500 ;
        RECT 90.830 161.810 91.000 162.500 ;
        RECT 91.420 161.810 91.590 162.500 ;
        RECT 92.330 161.810 92.500 162.500 ;
        RECT 92.920 161.810 93.090 162.500 ;
        RECT 93.830 161.810 94.000 162.500 ;
        RECT 94.420 161.810 94.590 162.500 ;
        RECT 95.330 161.810 95.500 162.500 ;
        RECT 84.210 161.470 84.710 161.640 ;
        RECT 85.710 161.470 86.210 161.640 ;
        RECT 87.210 161.470 87.710 161.640 ;
        RECT 88.710 161.470 89.210 161.640 ;
        RECT 90.210 161.470 90.710 161.640 ;
        RECT 91.710 161.470 92.210 161.640 ;
        RECT 93.210 161.470 93.710 161.640 ;
        RECT 94.710 161.470 95.210 161.640 ;
        RECT 95.990 161.175 96.160 163.135 ;
        RECT 83.210 161.005 96.160 161.175 ;
        RECT 42.920 159.955 55.620 160.125 ;
        RECT 42.920 157.645 43.090 159.955 ;
        RECT 43.770 159.535 44.270 159.705 ;
        RECT 45.270 159.535 45.770 159.705 ;
        RECT 46.770 159.535 47.270 159.705 ;
        RECT 48.270 159.535 48.770 159.705 ;
        RECT 49.770 159.535 50.270 159.705 ;
        RECT 51.270 159.535 51.770 159.705 ;
        RECT 52.770 159.535 53.270 159.705 ;
        RECT 54.270 159.535 54.770 159.705 ;
        RECT 43.480 158.280 43.650 159.320 ;
        RECT 44.390 158.280 44.560 159.320 ;
        RECT 44.980 158.280 45.150 159.320 ;
        RECT 45.890 158.280 46.060 159.320 ;
        RECT 46.480 158.280 46.650 159.320 ;
        RECT 47.390 158.280 47.560 159.320 ;
        RECT 47.980 158.280 48.150 159.320 ;
        RECT 48.890 158.280 49.060 159.320 ;
        RECT 49.480 158.280 49.650 159.320 ;
        RECT 50.390 158.280 50.560 159.320 ;
        RECT 50.980 158.280 51.150 159.320 ;
        RECT 51.890 158.280 52.060 159.320 ;
        RECT 52.480 158.280 52.650 159.320 ;
        RECT 53.390 158.280 53.560 159.320 ;
        RECT 53.980 158.280 54.150 159.320 ;
        RECT 54.890 158.280 55.060 159.320 ;
        RECT 43.770 157.895 44.270 158.065 ;
        RECT 45.270 157.895 45.770 158.065 ;
        RECT 46.770 157.895 47.270 158.065 ;
        RECT 48.270 157.895 48.770 158.065 ;
        RECT 49.770 157.895 50.270 158.065 ;
        RECT 51.270 157.895 51.770 158.065 ;
        RECT 52.770 157.895 53.270 158.065 ;
        RECT 54.270 157.895 54.770 158.065 ;
        RECT 55.450 157.645 55.620 159.955 ;
        RECT 42.920 157.475 55.620 157.645 ;
        RECT 56.400 159.955 69.100 160.125 ;
        RECT 56.400 157.645 56.570 159.955 ;
        RECT 57.250 159.535 57.750 159.705 ;
        RECT 58.750 159.535 59.250 159.705 ;
        RECT 60.250 159.535 60.750 159.705 ;
        RECT 61.750 159.535 62.250 159.705 ;
        RECT 63.250 159.535 63.750 159.705 ;
        RECT 64.750 159.535 65.250 159.705 ;
        RECT 66.250 159.535 66.750 159.705 ;
        RECT 67.750 159.535 68.250 159.705 ;
        RECT 56.960 158.280 57.130 159.320 ;
        RECT 57.870 158.280 58.040 159.320 ;
        RECT 58.460 158.280 58.630 159.320 ;
        RECT 59.370 158.280 59.540 159.320 ;
        RECT 59.960 158.280 60.130 159.320 ;
        RECT 60.870 158.280 61.040 159.320 ;
        RECT 61.460 158.280 61.630 159.320 ;
        RECT 62.370 158.280 62.540 159.320 ;
        RECT 62.960 158.280 63.130 159.320 ;
        RECT 63.870 158.280 64.040 159.320 ;
        RECT 64.460 158.280 64.630 159.320 ;
        RECT 65.370 158.280 65.540 159.320 ;
        RECT 65.960 158.280 66.130 159.320 ;
        RECT 66.870 158.280 67.040 159.320 ;
        RECT 67.460 158.280 67.630 159.320 ;
        RECT 68.370 158.280 68.540 159.320 ;
        RECT 57.250 157.895 57.750 158.065 ;
        RECT 58.750 157.895 59.250 158.065 ;
        RECT 60.250 157.895 60.750 158.065 ;
        RECT 61.750 157.895 62.250 158.065 ;
        RECT 63.250 157.895 63.750 158.065 ;
        RECT 64.750 157.895 65.250 158.065 ;
        RECT 66.250 157.895 66.750 158.065 ;
        RECT 67.750 157.895 68.250 158.065 ;
        RECT 68.930 157.645 69.100 159.955 ;
        RECT 56.400 157.475 69.100 157.645 ;
        RECT 69.880 159.955 82.580 160.125 ;
        RECT 69.880 157.645 70.050 159.955 ;
        RECT 70.730 159.535 71.230 159.705 ;
        RECT 72.230 159.535 72.730 159.705 ;
        RECT 73.730 159.535 74.230 159.705 ;
        RECT 75.230 159.535 75.730 159.705 ;
        RECT 76.730 159.535 77.230 159.705 ;
        RECT 78.230 159.535 78.730 159.705 ;
        RECT 79.730 159.535 80.230 159.705 ;
        RECT 81.230 159.535 81.730 159.705 ;
        RECT 70.440 158.280 70.610 159.320 ;
        RECT 71.350 158.280 71.520 159.320 ;
        RECT 71.940 158.280 72.110 159.320 ;
        RECT 72.850 158.280 73.020 159.320 ;
        RECT 73.440 158.280 73.610 159.320 ;
        RECT 74.350 158.280 74.520 159.320 ;
        RECT 74.940 158.280 75.110 159.320 ;
        RECT 75.850 158.280 76.020 159.320 ;
        RECT 76.440 158.280 76.610 159.320 ;
        RECT 77.350 158.280 77.520 159.320 ;
        RECT 77.940 158.280 78.110 159.320 ;
        RECT 78.850 158.280 79.020 159.320 ;
        RECT 79.440 158.280 79.610 159.320 ;
        RECT 80.350 158.280 80.520 159.320 ;
        RECT 80.940 158.280 81.110 159.320 ;
        RECT 81.850 158.280 82.020 159.320 ;
        RECT 70.730 157.895 71.230 158.065 ;
        RECT 72.230 157.895 72.730 158.065 ;
        RECT 73.730 157.895 74.230 158.065 ;
        RECT 75.230 157.895 75.730 158.065 ;
        RECT 76.730 157.895 77.230 158.065 ;
        RECT 78.230 157.895 78.730 158.065 ;
        RECT 79.730 157.895 80.230 158.065 ;
        RECT 81.230 157.895 81.730 158.065 ;
        RECT 82.410 157.645 82.580 159.955 ;
        RECT 69.880 157.475 82.580 157.645 ;
        RECT 83.360 159.955 96.060 160.125 ;
        RECT 83.360 157.645 83.530 159.955 ;
        RECT 84.210 159.535 84.710 159.705 ;
        RECT 85.710 159.535 86.210 159.705 ;
        RECT 87.210 159.535 87.710 159.705 ;
        RECT 88.710 159.535 89.210 159.705 ;
        RECT 90.210 159.535 90.710 159.705 ;
        RECT 91.710 159.535 92.210 159.705 ;
        RECT 93.210 159.535 93.710 159.705 ;
        RECT 94.710 159.535 95.210 159.705 ;
        RECT 83.920 158.280 84.090 159.320 ;
        RECT 84.830 158.280 85.000 159.320 ;
        RECT 85.420 158.280 85.590 159.320 ;
        RECT 86.330 158.280 86.500 159.320 ;
        RECT 86.920 158.280 87.090 159.320 ;
        RECT 87.830 158.280 88.000 159.320 ;
        RECT 88.420 158.280 88.590 159.320 ;
        RECT 89.330 158.280 89.500 159.320 ;
        RECT 89.920 158.280 90.090 159.320 ;
        RECT 90.830 158.280 91.000 159.320 ;
        RECT 91.420 158.280 91.590 159.320 ;
        RECT 92.330 158.280 92.500 159.320 ;
        RECT 92.920 158.280 93.090 159.320 ;
        RECT 93.830 158.280 94.000 159.320 ;
        RECT 94.420 158.280 94.590 159.320 ;
        RECT 95.330 158.280 95.500 159.320 ;
        RECT 84.210 157.895 84.710 158.065 ;
        RECT 85.710 157.895 86.210 158.065 ;
        RECT 87.210 157.895 87.710 158.065 ;
        RECT 88.710 157.895 89.210 158.065 ;
        RECT 90.210 157.895 90.710 158.065 ;
        RECT 91.710 157.895 92.210 158.065 ;
        RECT 93.210 157.895 93.710 158.065 ;
        RECT 94.710 157.895 95.210 158.065 ;
        RECT 95.890 157.645 96.060 159.955 ;
        RECT 83.360 157.475 96.060 157.645 ;
        RECT 36.205 154.605 38.505 154.775 ;
        RECT 36.205 140.495 36.375 154.605 ;
        RECT 37.010 153.945 37.700 154.115 ;
        RECT 36.670 153.325 36.840 153.825 ;
        RECT 37.870 153.325 38.040 153.825 ;
        RECT 37.010 153.035 37.700 153.205 ;
        RECT 37.010 152.445 37.700 152.615 ;
        RECT 36.670 151.825 36.840 152.325 ;
        RECT 37.870 151.825 38.040 152.325 ;
        RECT 37.010 151.535 37.700 151.705 ;
        RECT 37.010 150.945 37.700 151.115 ;
        RECT 36.670 150.325 36.840 150.825 ;
        RECT 37.870 150.325 38.040 150.825 ;
        RECT 37.010 150.035 37.700 150.205 ;
        RECT 37.010 149.445 37.700 149.615 ;
        RECT 36.670 148.825 36.840 149.325 ;
        RECT 37.870 148.825 38.040 149.325 ;
        RECT 37.010 148.535 37.700 148.705 ;
        RECT 37.010 147.945 37.700 148.115 ;
        RECT 36.670 147.325 36.840 147.825 ;
        RECT 37.870 147.325 38.040 147.825 ;
        RECT 37.010 147.035 37.700 147.205 ;
        RECT 37.010 146.445 37.700 146.615 ;
        RECT 36.670 145.825 36.840 146.325 ;
        RECT 37.870 145.825 38.040 146.325 ;
        RECT 37.010 145.535 37.700 145.705 ;
        RECT 37.010 144.945 37.700 145.115 ;
        RECT 36.670 144.325 36.840 144.825 ;
        RECT 37.870 144.325 38.040 144.825 ;
        RECT 37.010 144.035 37.700 144.205 ;
        RECT 37.010 143.445 37.700 143.615 ;
        RECT 36.670 142.825 36.840 143.325 ;
        RECT 37.870 142.825 38.040 143.325 ;
        RECT 37.010 142.535 37.700 142.705 ;
        RECT 37.010 141.945 37.700 142.115 ;
        RECT 36.670 141.325 36.840 141.825 ;
        RECT 37.870 141.325 38.040 141.825 ;
        RECT 37.010 141.035 37.700 141.205 ;
        RECT 38.335 140.495 38.505 154.605 ;
        RECT 36.205 140.325 38.505 140.495 ;
        RECT 39.385 154.505 42.035 154.675 ;
        RECT 39.385 140.645 39.555 154.505 ;
        RECT 40.190 153.945 41.230 154.115 ;
        RECT 39.805 153.325 39.975 153.825 ;
        RECT 41.445 153.325 41.615 153.825 ;
        RECT 40.190 153.035 41.230 153.205 ;
        RECT 40.190 152.445 41.230 152.615 ;
        RECT 39.805 151.825 39.975 152.325 ;
        RECT 41.445 151.825 41.615 152.325 ;
        RECT 40.190 151.535 41.230 151.705 ;
        RECT 40.190 150.945 41.230 151.115 ;
        RECT 39.805 150.325 39.975 150.825 ;
        RECT 41.445 150.325 41.615 150.825 ;
        RECT 40.190 150.035 41.230 150.205 ;
        RECT 40.190 149.445 41.230 149.615 ;
        RECT 39.805 148.825 39.975 149.325 ;
        RECT 41.445 148.825 41.615 149.325 ;
        RECT 40.190 148.535 41.230 148.705 ;
        RECT 40.190 147.945 41.230 148.115 ;
        RECT 39.805 147.325 39.975 147.825 ;
        RECT 41.445 147.325 41.615 147.825 ;
        RECT 40.190 147.035 41.230 147.205 ;
        RECT 40.190 146.445 41.230 146.615 ;
        RECT 39.805 145.825 39.975 146.325 ;
        RECT 41.445 145.825 41.615 146.325 ;
        RECT 40.190 145.535 41.230 145.705 ;
        RECT 40.190 144.945 41.230 145.115 ;
        RECT 39.805 144.325 39.975 144.825 ;
        RECT 41.445 144.325 41.615 144.825 ;
        RECT 40.190 144.035 41.230 144.205 ;
        RECT 40.190 143.445 41.230 143.615 ;
        RECT 39.805 142.825 39.975 143.325 ;
        RECT 41.445 142.825 41.615 143.325 ;
        RECT 40.190 142.535 41.230 142.705 ;
        RECT 40.190 141.945 41.230 142.115 ;
        RECT 39.805 141.325 39.975 141.825 ;
        RECT 41.445 141.325 41.615 141.825 ;
        RECT 40.190 141.035 41.230 141.205 ;
        RECT 41.865 140.645 42.035 154.505 ;
        RECT 39.385 140.475 42.035 140.645 ;
        RECT 42.915 154.605 45.215 154.775 ;
        RECT 42.915 140.495 43.085 154.605 ;
        RECT 43.720 153.945 44.410 154.115 ;
        RECT 43.380 153.325 43.550 153.825 ;
        RECT 44.580 153.325 44.750 153.825 ;
        RECT 43.720 153.035 44.410 153.205 ;
        RECT 43.720 152.445 44.410 152.615 ;
        RECT 43.380 151.825 43.550 152.325 ;
        RECT 44.580 151.825 44.750 152.325 ;
        RECT 43.720 151.535 44.410 151.705 ;
        RECT 43.720 150.945 44.410 151.115 ;
        RECT 43.380 150.325 43.550 150.825 ;
        RECT 44.580 150.325 44.750 150.825 ;
        RECT 43.720 150.035 44.410 150.205 ;
        RECT 43.720 149.445 44.410 149.615 ;
        RECT 43.380 148.825 43.550 149.325 ;
        RECT 44.580 148.825 44.750 149.325 ;
        RECT 43.720 148.535 44.410 148.705 ;
        RECT 43.720 147.945 44.410 148.115 ;
        RECT 43.380 147.325 43.550 147.825 ;
        RECT 44.580 147.325 44.750 147.825 ;
        RECT 43.720 147.035 44.410 147.205 ;
        RECT 43.720 146.445 44.410 146.615 ;
        RECT 43.380 145.825 43.550 146.325 ;
        RECT 44.580 145.825 44.750 146.325 ;
        RECT 43.720 145.535 44.410 145.705 ;
        RECT 43.720 144.945 44.410 145.115 ;
        RECT 43.380 144.325 43.550 144.825 ;
        RECT 44.580 144.325 44.750 144.825 ;
        RECT 43.720 144.035 44.410 144.205 ;
        RECT 43.720 143.445 44.410 143.615 ;
        RECT 43.380 142.825 43.550 143.325 ;
        RECT 44.580 142.825 44.750 143.325 ;
        RECT 43.720 142.535 44.410 142.705 ;
        RECT 43.720 141.945 44.410 142.115 ;
        RECT 43.380 141.325 43.550 141.825 ;
        RECT 44.580 141.325 44.750 141.825 ;
        RECT 43.720 141.035 44.410 141.205 ;
        RECT 45.045 140.495 45.215 154.605 ;
        RECT 42.915 140.325 45.215 140.495 ;
        RECT 46.095 154.505 48.745 154.675 ;
        RECT 46.095 140.645 46.265 154.505 ;
        RECT 46.900 153.945 47.940 154.115 ;
        RECT 46.515 153.325 46.685 153.825 ;
        RECT 48.155 153.325 48.325 153.825 ;
        RECT 46.900 153.035 47.940 153.205 ;
        RECT 46.900 152.445 47.940 152.615 ;
        RECT 46.515 151.825 46.685 152.325 ;
        RECT 48.155 151.825 48.325 152.325 ;
        RECT 46.900 151.535 47.940 151.705 ;
        RECT 46.900 150.945 47.940 151.115 ;
        RECT 46.515 150.325 46.685 150.825 ;
        RECT 48.155 150.325 48.325 150.825 ;
        RECT 46.900 150.035 47.940 150.205 ;
        RECT 46.900 149.445 47.940 149.615 ;
        RECT 46.515 148.825 46.685 149.325 ;
        RECT 48.155 148.825 48.325 149.325 ;
        RECT 46.900 148.535 47.940 148.705 ;
        RECT 46.900 147.945 47.940 148.115 ;
        RECT 46.515 147.325 46.685 147.825 ;
        RECT 48.155 147.325 48.325 147.825 ;
        RECT 46.900 147.035 47.940 147.205 ;
        RECT 46.900 146.445 47.940 146.615 ;
        RECT 46.515 145.825 46.685 146.325 ;
        RECT 48.155 145.825 48.325 146.325 ;
        RECT 46.900 145.535 47.940 145.705 ;
        RECT 46.900 144.945 47.940 145.115 ;
        RECT 46.515 144.325 46.685 144.825 ;
        RECT 48.155 144.325 48.325 144.825 ;
        RECT 46.900 144.035 47.940 144.205 ;
        RECT 46.900 143.445 47.940 143.615 ;
        RECT 46.515 142.825 46.685 143.325 ;
        RECT 48.155 142.825 48.325 143.325 ;
        RECT 46.900 142.535 47.940 142.705 ;
        RECT 46.900 141.945 47.940 142.115 ;
        RECT 46.515 141.325 46.685 141.825 ;
        RECT 48.155 141.325 48.325 141.825 ;
        RECT 46.900 141.035 47.940 141.205 ;
        RECT 48.575 140.645 48.745 154.505 ;
        RECT 46.095 140.475 48.745 140.645 ;
        RECT 49.625 154.605 51.925 154.775 ;
        RECT 49.625 140.495 49.795 154.605 ;
        RECT 50.430 153.945 51.120 154.115 ;
        RECT 50.090 153.325 50.260 153.825 ;
        RECT 51.290 153.325 51.460 153.825 ;
        RECT 50.430 153.035 51.120 153.205 ;
        RECT 50.430 152.445 51.120 152.615 ;
        RECT 50.090 151.825 50.260 152.325 ;
        RECT 51.290 151.825 51.460 152.325 ;
        RECT 50.430 151.535 51.120 151.705 ;
        RECT 50.430 150.945 51.120 151.115 ;
        RECT 50.090 150.325 50.260 150.825 ;
        RECT 51.290 150.325 51.460 150.825 ;
        RECT 50.430 150.035 51.120 150.205 ;
        RECT 50.430 149.445 51.120 149.615 ;
        RECT 50.090 148.825 50.260 149.325 ;
        RECT 51.290 148.825 51.460 149.325 ;
        RECT 50.430 148.535 51.120 148.705 ;
        RECT 50.430 147.945 51.120 148.115 ;
        RECT 50.090 147.325 50.260 147.825 ;
        RECT 51.290 147.325 51.460 147.825 ;
        RECT 50.430 147.035 51.120 147.205 ;
        RECT 50.430 146.445 51.120 146.615 ;
        RECT 50.090 145.825 50.260 146.325 ;
        RECT 51.290 145.825 51.460 146.325 ;
        RECT 50.430 145.535 51.120 145.705 ;
        RECT 50.430 144.945 51.120 145.115 ;
        RECT 50.090 144.325 50.260 144.825 ;
        RECT 51.290 144.325 51.460 144.825 ;
        RECT 50.430 144.035 51.120 144.205 ;
        RECT 50.430 143.445 51.120 143.615 ;
        RECT 50.090 142.825 50.260 143.325 ;
        RECT 51.290 142.825 51.460 143.325 ;
        RECT 50.430 142.535 51.120 142.705 ;
        RECT 50.430 141.945 51.120 142.115 ;
        RECT 50.090 141.325 50.260 141.825 ;
        RECT 51.290 141.325 51.460 141.825 ;
        RECT 50.430 141.035 51.120 141.205 ;
        RECT 51.755 140.495 51.925 154.605 ;
        RECT 49.625 140.325 51.925 140.495 ;
        RECT 52.805 154.505 55.455 154.675 ;
        RECT 52.805 140.645 52.975 154.505 ;
        RECT 53.610 153.945 54.650 154.115 ;
        RECT 53.225 153.325 53.395 153.825 ;
        RECT 54.865 153.325 55.035 153.825 ;
        RECT 53.610 153.035 54.650 153.205 ;
        RECT 53.610 152.445 54.650 152.615 ;
        RECT 53.225 151.825 53.395 152.325 ;
        RECT 54.865 151.825 55.035 152.325 ;
        RECT 53.610 151.535 54.650 151.705 ;
        RECT 53.610 150.945 54.650 151.115 ;
        RECT 53.225 150.325 53.395 150.825 ;
        RECT 54.865 150.325 55.035 150.825 ;
        RECT 53.610 150.035 54.650 150.205 ;
        RECT 53.610 149.445 54.650 149.615 ;
        RECT 53.225 148.825 53.395 149.325 ;
        RECT 54.865 148.825 55.035 149.325 ;
        RECT 53.610 148.535 54.650 148.705 ;
        RECT 53.610 147.945 54.650 148.115 ;
        RECT 53.225 147.325 53.395 147.825 ;
        RECT 54.865 147.325 55.035 147.825 ;
        RECT 53.610 147.035 54.650 147.205 ;
        RECT 53.610 146.445 54.650 146.615 ;
        RECT 53.225 145.825 53.395 146.325 ;
        RECT 54.865 145.825 55.035 146.325 ;
        RECT 53.610 145.535 54.650 145.705 ;
        RECT 53.610 144.945 54.650 145.115 ;
        RECT 53.225 144.325 53.395 144.825 ;
        RECT 54.865 144.325 55.035 144.825 ;
        RECT 53.610 144.035 54.650 144.205 ;
        RECT 53.610 143.445 54.650 143.615 ;
        RECT 53.225 142.825 53.395 143.325 ;
        RECT 54.865 142.825 55.035 143.325 ;
        RECT 53.610 142.535 54.650 142.705 ;
        RECT 53.610 141.945 54.650 142.115 ;
        RECT 53.225 141.325 53.395 141.825 ;
        RECT 54.865 141.325 55.035 141.825 ;
        RECT 53.610 141.035 54.650 141.205 ;
        RECT 55.285 140.645 55.455 154.505 ;
        RECT 52.805 140.475 55.455 140.645 ;
        RECT 56.335 154.605 58.635 154.775 ;
        RECT 56.335 140.495 56.505 154.605 ;
        RECT 57.140 153.945 57.830 154.115 ;
        RECT 56.800 153.325 56.970 153.825 ;
        RECT 58.000 153.325 58.170 153.825 ;
        RECT 57.140 153.035 57.830 153.205 ;
        RECT 57.140 152.445 57.830 152.615 ;
        RECT 56.800 151.825 56.970 152.325 ;
        RECT 58.000 151.825 58.170 152.325 ;
        RECT 57.140 151.535 57.830 151.705 ;
        RECT 57.140 150.945 57.830 151.115 ;
        RECT 56.800 150.325 56.970 150.825 ;
        RECT 58.000 150.325 58.170 150.825 ;
        RECT 57.140 150.035 57.830 150.205 ;
        RECT 57.140 149.445 57.830 149.615 ;
        RECT 56.800 148.825 56.970 149.325 ;
        RECT 58.000 148.825 58.170 149.325 ;
        RECT 57.140 148.535 57.830 148.705 ;
        RECT 57.140 147.945 57.830 148.115 ;
        RECT 56.800 147.325 56.970 147.825 ;
        RECT 58.000 147.325 58.170 147.825 ;
        RECT 57.140 147.035 57.830 147.205 ;
        RECT 57.140 146.445 57.830 146.615 ;
        RECT 56.800 145.825 56.970 146.325 ;
        RECT 58.000 145.825 58.170 146.325 ;
        RECT 57.140 145.535 57.830 145.705 ;
        RECT 57.140 144.945 57.830 145.115 ;
        RECT 56.800 144.325 56.970 144.825 ;
        RECT 58.000 144.325 58.170 144.825 ;
        RECT 57.140 144.035 57.830 144.205 ;
        RECT 57.140 143.445 57.830 143.615 ;
        RECT 56.800 142.825 56.970 143.325 ;
        RECT 58.000 142.825 58.170 143.325 ;
        RECT 57.140 142.535 57.830 142.705 ;
        RECT 57.140 141.945 57.830 142.115 ;
        RECT 56.800 141.325 56.970 141.825 ;
        RECT 58.000 141.325 58.170 141.825 ;
        RECT 57.140 141.035 57.830 141.205 ;
        RECT 58.465 140.495 58.635 154.605 ;
        RECT 56.335 140.325 58.635 140.495 ;
        RECT 59.515 154.505 62.165 154.675 ;
        RECT 59.515 140.645 59.685 154.505 ;
        RECT 60.320 153.945 61.360 154.115 ;
        RECT 59.935 153.325 60.105 153.825 ;
        RECT 61.575 153.325 61.745 153.825 ;
        RECT 60.320 153.035 61.360 153.205 ;
        RECT 60.320 152.445 61.360 152.615 ;
        RECT 59.935 151.825 60.105 152.325 ;
        RECT 61.575 151.825 61.745 152.325 ;
        RECT 60.320 151.535 61.360 151.705 ;
        RECT 60.320 150.945 61.360 151.115 ;
        RECT 59.935 150.325 60.105 150.825 ;
        RECT 61.575 150.325 61.745 150.825 ;
        RECT 60.320 150.035 61.360 150.205 ;
        RECT 60.320 149.445 61.360 149.615 ;
        RECT 59.935 148.825 60.105 149.325 ;
        RECT 61.575 148.825 61.745 149.325 ;
        RECT 60.320 148.535 61.360 148.705 ;
        RECT 60.320 147.945 61.360 148.115 ;
        RECT 59.935 147.325 60.105 147.825 ;
        RECT 61.575 147.325 61.745 147.825 ;
        RECT 60.320 147.035 61.360 147.205 ;
        RECT 60.320 146.445 61.360 146.615 ;
        RECT 59.935 145.825 60.105 146.325 ;
        RECT 61.575 145.825 61.745 146.325 ;
        RECT 60.320 145.535 61.360 145.705 ;
        RECT 60.320 144.945 61.360 145.115 ;
        RECT 59.935 144.325 60.105 144.825 ;
        RECT 61.575 144.325 61.745 144.825 ;
        RECT 60.320 144.035 61.360 144.205 ;
        RECT 60.320 143.445 61.360 143.615 ;
        RECT 59.935 142.825 60.105 143.325 ;
        RECT 61.575 142.825 61.745 143.325 ;
        RECT 60.320 142.535 61.360 142.705 ;
        RECT 60.320 141.945 61.360 142.115 ;
        RECT 59.935 141.325 60.105 141.825 ;
        RECT 61.575 141.325 61.745 141.825 ;
        RECT 60.320 141.035 61.360 141.205 ;
        RECT 61.995 140.645 62.165 154.505 ;
        RECT 59.515 140.475 62.165 140.645 ;
        RECT 63.045 154.605 65.345 154.775 ;
        RECT 63.045 140.495 63.215 154.605 ;
        RECT 63.850 153.945 64.540 154.115 ;
        RECT 63.510 153.325 63.680 153.825 ;
        RECT 64.710 153.325 64.880 153.825 ;
        RECT 63.850 153.035 64.540 153.205 ;
        RECT 63.850 152.445 64.540 152.615 ;
        RECT 63.510 151.825 63.680 152.325 ;
        RECT 64.710 151.825 64.880 152.325 ;
        RECT 63.850 151.535 64.540 151.705 ;
        RECT 63.850 150.945 64.540 151.115 ;
        RECT 63.510 150.325 63.680 150.825 ;
        RECT 64.710 150.325 64.880 150.825 ;
        RECT 63.850 150.035 64.540 150.205 ;
        RECT 63.850 149.445 64.540 149.615 ;
        RECT 63.510 148.825 63.680 149.325 ;
        RECT 64.710 148.825 64.880 149.325 ;
        RECT 63.850 148.535 64.540 148.705 ;
        RECT 63.850 147.945 64.540 148.115 ;
        RECT 63.510 147.325 63.680 147.825 ;
        RECT 64.710 147.325 64.880 147.825 ;
        RECT 63.850 147.035 64.540 147.205 ;
        RECT 63.850 146.445 64.540 146.615 ;
        RECT 63.510 145.825 63.680 146.325 ;
        RECT 64.710 145.825 64.880 146.325 ;
        RECT 63.850 145.535 64.540 145.705 ;
        RECT 63.850 144.945 64.540 145.115 ;
        RECT 63.510 144.325 63.680 144.825 ;
        RECT 64.710 144.325 64.880 144.825 ;
        RECT 63.850 144.035 64.540 144.205 ;
        RECT 63.850 143.445 64.540 143.615 ;
        RECT 63.510 142.825 63.680 143.325 ;
        RECT 64.710 142.825 64.880 143.325 ;
        RECT 63.850 142.535 64.540 142.705 ;
        RECT 63.850 141.945 64.540 142.115 ;
        RECT 63.510 141.325 63.680 141.825 ;
        RECT 64.710 141.325 64.880 141.825 ;
        RECT 63.850 141.035 64.540 141.205 ;
        RECT 65.175 140.495 65.345 154.605 ;
        RECT 63.045 140.325 65.345 140.495 ;
        RECT 66.225 154.505 68.875 154.675 ;
        RECT 66.225 140.645 66.395 154.505 ;
        RECT 67.030 153.945 68.070 154.115 ;
        RECT 66.645 153.325 66.815 153.825 ;
        RECT 68.285 153.325 68.455 153.825 ;
        RECT 67.030 153.035 68.070 153.205 ;
        RECT 67.030 152.445 68.070 152.615 ;
        RECT 66.645 151.825 66.815 152.325 ;
        RECT 68.285 151.825 68.455 152.325 ;
        RECT 67.030 151.535 68.070 151.705 ;
        RECT 67.030 150.945 68.070 151.115 ;
        RECT 66.645 150.325 66.815 150.825 ;
        RECT 68.285 150.325 68.455 150.825 ;
        RECT 67.030 150.035 68.070 150.205 ;
        RECT 67.030 149.445 68.070 149.615 ;
        RECT 66.645 148.825 66.815 149.325 ;
        RECT 68.285 148.825 68.455 149.325 ;
        RECT 67.030 148.535 68.070 148.705 ;
        RECT 67.030 147.945 68.070 148.115 ;
        RECT 66.645 147.325 66.815 147.825 ;
        RECT 68.285 147.325 68.455 147.825 ;
        RECT 67.030 147.035 68.070 147.205 ;
        RECT 67.030 146.445 68.070 146.615 ;
        RECT 66.645 145.825 66.815 146.325 ;
        RECT 68.285 145.825 68.455 146.325 ;
        RECT 67.030 145.535 68.070 145.705 ;
        RECT 67.030 144.945 68.070 145.115 ;
        RECT 66.645 144.325 66.815 144.825 ;
        RECT 68.285 144.325 68.455 144.825 ;
        RECT 67.030 144.035 68.070 144.205 ;
        RECT 67.030 143.445 68.070 143.615 ;
        RECT 66.645 142.825 66.815 143.325 ;
        RECT 68.285 142.825 68.455 143.325 ;
        RECT 67.030 142.535 68.070 142.705 ;
        RECT 67.030 141.945 68.070 142.115 ;
        RECT 66.645 141.325 66.815 141.825 ;
        RECT 68.285 141.325 68.455 141.825 ;
        RECT 67.030 141.035 68.070 141.205 ;
        RECT 68.705 140.645 68.875 154.505 ;
        RECT 66.225 140.475 68.875 140.645 ;
        RECT 69.755 154.605 72.055 154.775 ;
        RECT 69.755 140.495 69.925 154.605 ;
        RECT 70.560 153.945 71.250 154.115 ;
        RECT 70.220 153.325 70.390 153.825 ;
        RECT 71.420 153.325 71.590 153.825 ;
        RECT 70.560 153.035 71.250 153.205 ;
        RECT 70.560 152.445 71.250 152.615 ;
        RECT 70.220 151.825 70.390 152.325 ;
        RECT 71.420 151.825 71.590 152.325 ;
        RECT 70.560 151.535 71.250 151.705 ;
        RECT 70.560 150.945 71.250 151.115 ;
        RECT 70.220 150.325 70.390 150.825 ;
        RECT 71.420 150.325 71.590 150.825 ;
        RECT 70.560 150.035 71.250 150.205 ;
        RECT 70.560 149.445 71.250 149.615 ;
        RECT 70.220 148.825 70.390 149.325 ;
        RECT 71.420 148.825 71.590 149.325 ;
        RECT 70.560 148.535 71.250 148.705 ;
        RECT 70.560 147.945 71.250 148.115 ;
        RECT 70.220 147.325 70.390 147.825 ;
        RECT 71.420 147.325 71.590 147.825 ;
        RECT 70.560 147.035 71.250 147.205 ;
        RECT 70.560 146.445 71.250 146.615 ;
        RECT 70.220 145.825 70.390 146.325 ;
        RECT 71.420 145.825 71.590 146.325 ;
        RECT 70.560 145.535 71.250 145.705 ;
        RECT 70.560 144.945 71.250 145.115 ;
        RECT 70.220 144.325 70.390 144.825 ;
        RECT 71.420 144.325 71.590 144.825 ;
        RECT 70.560 144.035 71.250 144.205 ;
        RECT 70.560 143.445 71.250 143.615 ;
        RECT 70.220 142.825 70.390 143.325 ;
        RECT 71.420 142.825 71.590 143.325 ;
        RECT 70.560 142.535 71.250 142.705 ;
        RECT 70.560 141.945 71.250 142.115 ;
        RECT 70.220 141.325 70.390 141.825 ;
        RECT 71.420 141.325 71.590 141.825 ;
        RECT 70.560 141.035 71.250 141.205 ;
        RECT 71.885 140.495 72.055 154.605 ;
        RECT 69.755 140.325 72.055 140.495 ;
        RECT 72.935 154.505 75.585 154.675 ;
        RECT 72.935 140.645 73.105 154.505 ;
        RECT 73.740 153.945 74.780 154.115 ;
        RECT 73.355 153.325 73.525 153.825 ;
        RECT 74.995 153.325 75.165 153.825 ;
        RECT 73.740 153.035 74.780 153.205 ;
        RECT 73.740 152.445 74.780 152.615 ;
        RECT 73.355 151.825 73.525 152.325 ;
        RECT 74.995 151.825 75.165 152.325 ;
        RECT 73.740 151.535 74.780 151.705 ;
        RECT 73.740 150.945 74.780 151.115 ;
        RECT 73.355 150.325 73.525 150.825 ;
        RECT 74.995 150.325 75.165 150.825 ;
        RECT 73.740 150.035 74.780 150.205 ;
        RECT 73.740 149.445 74.780 149.615 ;
        RECT 73.355 148.825 73.525 149.325 ;
        RECT 74.995 148.825 75.165 149.325 ;
        RECT 73.740 148.535 74.780 148.705 ;
        RECT 73.740 147.945 74.780 148.115 ;
        RECT 73.355 147.325 73.525 147.825 ;
        RECT 74.995 147.325 75.165 147.825 ;
        RECT 73.740 147.035 74.780 147.205 ;
        RECT 73.740 146.445 74.780 146.615 ;
        RECT 73.355 145.825 73.525 146.325 ;
        RECT 74.995 145.825 75.165 146.325 ;
        RECT 73.740 145.535 74.780 145.705 ;
        RECT 73.740 144.945 74.780 145.115 ;
        RECT 73.355 144.325 73.525 144.825 ;
        RECT 74.995 144.325 75.165 144.825 ;
        RECT 73.740 144.035 74.780 144.205 ;
        RECT 73.740 143.445 74.780 143.615 ;
        RECT 73.355 142.825 73.525 143.325 ;
        RECT 74.995 142.825 75.165 143.325 ;
        RECT 73.740 142.535 74.780 142.705 ;
        RECT 73.740 141.945 74.780 142.115 ;
        RECT 73.355 141.325 73.525 141.825 ;
        RECT 74.995 141.325 75.165 141.825 ;
        RECT 73.740 141.035 74.780 141.205 ;
        RECT 75.415 140.645 75.585 154.505 ;
        RECT 72.935 140.475 75.585 140.645 ;
        RECT 76.465 154.605 78.765 154.775 ;
        RECT 76.465 140.495 76.635 154.605 ;
        RECT 77.270 153.945 77.960 154.115 ;
        RECT 76.930 153.325 77.100 153.825 ;
        RECT 78.130 153.325 78.300 153.825 ;
        RECT 77.270 153.035 77.960 153.205 ;
        RECT 77.270 152.445 77.960 152.615 ;
        RECT 76.930 151.825 77.100 152.325 ;
        RECT 78.130 151.825 78.300 152.325 ;
        RECT 77.270 151.535 77.960 151.705 ;
        RECT 77.270 150.945 77.960 151.115 ;
        RECT 76.930 150.325 77.100 150.825 ;
        RECT 78.130 150.325 78.300 150.825 ;
        RECT 77.270 150.035 77.960 150.205 ;
        RECT 77.270 149.445 77.960 149.615 ;
        RECT 76.930 148.825 77.100 149.325 ;
        RECT 78.130 148.825 78.300 149.325 ;
        RECT 77.270 148.535 77.960 148.705 ;
        RECT 77.270 147.945 77.960 148.115 ;
        RECT 76.930 147.325 77.100 147.825 ;
        RECT 78.130 147.325 78.300 147.825 ;
        RECT 77.270 147.035 77.960 147.205 ;
        RECT 77.270 146.445 77.960 146.615 ;
        RECT 76.930 145.825 77.100 146.325 ;
        RECT 78.130 145.825 78.300 146.325 ;
        RECT 77.270 145.535 77.960 145.705 ;
        RECT 77.270 144.945 77.960 145.115 ;
        RECT 76.930 144.325 77.100 144.825 ;
        RECT 78.130 144.325 78.300 144.825 ;
        RECT 77.270 144.035 77.960 144.205 ;
        RECT 77.270 143.445 77.960 143.615 ;
        RECT 76.930 142.825 77.100 143.325 ;
        RECT 78.130 142.825 78.300 143.325 ;
        RECT 77.270 142.535 77.960 142.705 ;
        RECT 77.270 141.945 77.960 142.115 ;
        RECT 76.930 141.325 77.100 141.825 ;
        RECT 78.130 141.325 78.300 141.825 ;
        RECT 77.270 141.035 77.960 141.205 ;
        RECT 78.595 140.495 78.765 154.605 ;
        RECT 76.465 140.325 78.765 140.495 ;
        RECT 79.645 154.505 82.295 154.675 ;
        RECT 79.645 140.645 79.815 154.505 ;
        RECT 80.450 153.945 81.490 154.115 ;
        RECT 80.065 153.325 80.235 153.825 ;
        RECT 81.705 153.325 81.875 153.825 ;
        RECT 80.450 153.035 81.490 153.205 ;
        RECT 80.450 152.445 81.490 152.615 ;
        RECT 80.065 151.825 80.235 152.325 ;
        RECT 81.705 151.825 81.875 152.325 ;
        RECT 80.450 151.535 81.490 151.705 ;
        RECT 80.450 150.945 81.490 151.115 ;
        RECT 80.065 150.325 80.235 150.825 ;
        RECT 81.705 150.325 81.875 150.825 ;
        RECT 80.450 150.035 81.490 150.205 ;
        RECT 80.450 149.445 81.490 149.615 ;
        RECT 80.065 148.825 80.235 149.325 ;
        RECT 81.705 148.825 81.875 149.325 ;
        RECT 80.450 148.535 81.490 148.705 ;
        RECT 80.450 147.945 81.490 148.115 ;
        RECT 80.065 147.325 80.235 147.825 ;
        RECT 81.705 147.325 81.875 147.825 ;
        RECT 80.450 147.035 81.490 147.205 ;
        RECT 80.450 146.445 81.490 146.615 ;
        RECT 80.065 145.825 80.235 146.325 ;
        RECT 81.705 145.825 81.875 146.325 ;
        RECT 80.450 145.535 81.490 145.705 ;
        RECT 80.450 144.945 81.490 145.115 ;
        RECT 80.065 144.325 80.235 144.825 ;
        RECT 81.705 144.325 81.875 144.825 ;
        RECT 80.450 144.035 81.490 144.205 ;
        RECT 80.450 143.445 81.490 143.615 ;
        RECT 80.065 142.825 80.235 143.325 ;
        RECT 81.705 142.825 81.875 143.325 ;
        RECT 80.450 142.535 81.490 142.705 ;
        RECT 80.450 141.945 81.490 142.115 ;
        RECT 80.065 141.325 80.235 141.825 ;
        RECT 81.705 141.325 81.875 141.825 ;
        RECT 80.450 141.035 81.490 141.205 ;
        RECT 82.125 140.645 82.295 154.505 ;
        RECT 79.645 140.475 82.295 140.645 ;
        RECT 83.175 154.605 85.475 154.775 ;
        RECT 83.175 140.495 83.345 154.605 ;
        RECT 83.980 153.945 84.670 154.115 ;
        RECT 83.640 153.325 83.810 153.825 ;
        RECT 84.840 153.325 85.010 153.825 ;
        RECT 83.980 153.035 84.670 153.205 ;
        RECT 83.980 152.445 84.670 152.615 ;
        RECT 83.640 151.825 83.810 152.325 ;
        RECT 84.840 151.825 85.010 152.325 ;
        RECT 83.980 151.535 84.670 151.705 ;
        RECT 83.980 150.945 84.670 151.115 ;
        RECT 83.640 150.325 83.810 150.825 ;
        RECT 84.840 150.325 85.010 150.825 ;
        RECT 83.980 150.035 84.670 150.205 ;
        RECT 83.980 149.445 84.670 149.615 ;
        RECT 83.640 148.825 83.810 149.325 ;
        RECT 84.840 148.825 85.010 149.325 ;
        RECT 83.980 148.535 84.670 148.705 ;
        RECT 83.980 147.945 84.670 148.115 ;
        RECT 83.640 147.325 83.810 147.825 ;
        RECT 84.840 147.325 85.010 147.825 ;
        RECT 83.980 147.035 84.670 147.205 ;
        RECT 83.980 146.445 84.670 146.615 ;
        RECT 83.640 145.825 83.810 146.325 ;
        RECT 84.840 145.825 85.010 146.325 ;
        RECT 83.980 145.535 84.670 145.705 ;
        RECT 83.980 144.945 84.670 145.115 ;
        RECT 83.640 144.325 83.810 144.825 ;
        RECT 84.840 144.325 85.010 144.825 ;
        RECT 83.980 144.035 84.670 144.205 ;
        RECT 83.980 143.445 84.670 143.615 ;
        RECT 83.640 142.825 83.810 143.325 ;
        RECT 84.840 142.825 85.010 143.325 ;
        RECT 83.980 142.535 84.670 142.705 ;
        RECT 83.980 141.945 84.670 142.115 ;
        RECT 83.640 141.325 83.810 141.825 ;
        RECT 84.840 141.325 85.010 141.825 ;
        RECT 83.980 141.035 84.670 141.205 ;
        RECT 85.305 140.495 85.475 154.605 ;
        RECT 83.175 140.325 85.475 140.495 ;
        RECT 86.355 154.505 89.005 154.675 ;
        RECT 86.355 140.645 86.525 154.505 ;
        RECT 87.160 153.945 88.200 154.115 ;
        RECT 86.775 153.325 86.945 153.825 ;
        RECT 88.415 153.325 88.585 153.825 ;
        RECT 87.160 153.035 88.200 153.205 ;
        RECT 87.160 152.445 88.200 152.615 ;
        RECT 86.775 151.825 86.945 152.325 ;
        RECT 88.415 151.825 88.585 152.325 ;
        RECT 87.160 151.535 88.200 151.705 ;
        RECT 87.160 150.945 88.200 151.115 ;
        RECT 86.775 150.325 86.945 150.825 ;
        RECT 88.415 150.325 88.585 150.825 ;
        RECT 87.160 150.035 88.200 150.205 ;
        RECT 87.160 149.445 88.200 149.615 ;
        RECT 86.775 148.825 86.945 149.325 ;
        RECT 88.415 148.825 88.585 149.325 ;
        RECT 87.160 148.535 88.200 148.705 ;
        RECT 87.160 147.945 88.200 148.115 ;
        RECT 86.775 147.325 86.945 147.825 ;
        RECT 88.415 147.325 88.585 147.825 ;
        RECT 87.160 147.035 88.200 147.205 ;
        RECT 87.160 146.445 88.200 146.615 ;
        RECT 86.775 145.825 86.945 146.325 ;
        RECT 88.415 145.825 88.585 146.325 ;
        RECT 87.160 145.535 88.200 145.705 ;
        RECT 87.160 144.945 88.200 145.115 ;
        RECT 86.775 144.325 86.945 144.825 ;
        RECT 88.415 144.325 88.585 144.825 ;
        RECT 87.160 144.035 88.200 144.205 ;
        RECT 87.160 143.445 88.200 143.615 ;
        RECT 86.775 142.825 86.945 143.325 ;
        RECT 88.415 142.825 88.585 143.325 ;
        RECT 87.160 142.535 88.200 142.705 ;
        RECT 87.160 141.945 88.200 142.115 ;
        RECT 86.775 141.325 86.945 141.825 ;
        RECT 88.415 141.325 88.585 141.825 ;
        RECT 87.160 141.035 88.200 141.205 ;
        RECT 88.835 140.645 89.005 154.505 ;
        RECT 86.355 140.475 89.005 140.645 ;
        RECT 89.885 154.605 92.185 154.775 ;
        RECT 89.885 140.495 90.055 154.605 ;
        RECT 90.690 153.945 91.380 154.115 ;
        RECT 90.350 153.325 90.520 153.825 ;
        RECT 91.550 153.325 91.720 153.825 ;
        RECT 90.690 153.035 91.380 153.205 ;
        RECT 90.690 152.445 91.380 152.615 ;
        RECT 90.350 151.825 90.520 152.325 ;
        RECT 91.550 151.825 91.720 152.325 ;
        RECT 90.690 151.535 91.380 151.705 ;
        RECT 90.690 150.945 91.380 151.115 ;
        RECT 90.350 150.325 90.520 150.825 ;
        RECT 91.550 150.325 91.720 150.825 ;
        RECT 90.690 150.035 91.380 150.205 ;
        RECT 90.690 149.445 91.380 149.615 ;
        RECT 90.350 148.825 90.520 149.325 ;
        RECT 91.550 148.825 91.720 149.325 ;
        RECT 90.690 148.535 91.380 148.705 ;
        RECT 90.690 147.945 91.380 148.115 ;
        RECT 90.350 147.325 90.520 147.825 ;
        RECT 91.550 147.325 91.720 147.825 ;
        RECT 90.690 147.035 91.380 147.205 ;
        RECT 90.690 146.445 91.380 146.615 ;
        RECT 90.350 145.825 90.520 146.325 ;
        RECT 91.550 145.825 91.720 146.325 ;
        RECT 90.690 145.535 91.380 145.705 ;
        RECT 90.690 144.945 91.380 145.115 ;
        RECT 90.350 144.325 90.520 144.825 ;
        RECT 91.550 144.325 91.720 144.825 ;
        RECT 90.690 144.035 91.380 144.205 ;
        RECT 90.690 143.445 91.380 143.615 ;
        RECT 90.350 142.825 90.520 143.325 ;
        RECT 91.550 142.825 91.720 143.325 ;
        RECT 90.690 142.535 91.380 142.705 ;
        RECT 90.690 141.945 91.380 142.115 ;
        RECT 90.350 141.325 90.520 141.825 ;
        RECT 91.550 141.325 91.720 141.825 ;
        RECT 90.690 141.035 91.380 141.205 ;
        RECT 92.015 140.495 92.185 154.605 ;
        RECT 89.885 140.325 92.185 140.495 ;
        RECT 93.065 154.505 95.715 154.675 ;
        RECT 93.065 140.645 93.235 154.505 ;
        RECT 93.870 153.945 94.910 154.115 ;
        RECT 93.485 153.325 93.655 153.825 ;
        RECT 95.125 153.325 95.295 153.825 ;
        RECT 93.870 153.035 94.910 153.205 ;
        RECT 93.870 152.445 94.910 152.615 ;
        RECT 93.485 151.825 93.655 152.325 ;
        RECT 95.125 151.825 95.295 152.325 ;
        RECT 93.870 151.535 94.910 151.705 ;
        RECT 93.870 150.945 94.910 151.115 ;
        RECT 93.485 150.325 93.655 150.825 ;
        RECT 95.125 150.325 95.295 150.825 ;
        RECT 93.870 150.035 94.910 150.205 ;
        RECT 93.870 149.445 94.910 149.615 ;
        RECT 93.485 148.825 93.655 149.325 ;
        RECT 95.125 148.825 95.295 149.325 ;
        RECT 93.870 148.535 94.910 148.705 ;
        RECT 93.870 147.945 94.910 148.115 ;
        RECT 93.485 147.325 93.655 147.825 ;
        RECT 95.125 147.325 95.295 147.825 ;
        RECT 93.870 147.035 94.910 147.205 ;
        RECT 93.870 146.445 94.910 146.615 ;
        RECT 93.485 145.825 93.655 146.325 ;
        RECT 95.125 145.825 95.295 146.325 ;
        RECT 93.870 145.535 94.910 145.705 ;
        RECT 93.870 144.945 94.910 145.115 ;
        RECT 93.485 144.325 93.655 144.825 ;
        RECT 95.125 144.325 95.295 144.825 ;
        RECT 93.870 144.035 94.910 144.205 ;
        RECT 93.870 143.445 94.910 143.615 ;
        RECT 93.485 142.825 93.655 143.325 ;
        RECT 95.125 142.825 95.295 143.325 ;
        RECT 93.870 142.535 94.910 142.705 ;
        RECT 93.870 141.945 94.910 142.115 ;
        RECT 93.485 141.325 93.655 141.825 ;
        RECT 95.125 141.325 95.295 141.825 ;
        RECT 93.870 141.035 94.910 141.205 ;
        RECT 95.545 140.645 95.715 154.505 ;
        RECT 93.065 140.475 95.715 140.645 ;
        RECT 96.595 154.605 98.895 154.775 ;
        RECT 96.595 140.495 96.765 154.605 ;
        RECT 97.400 153.945 98.090 154.115 ;
        RECT 97.060 153.325 97.230 153.825 ;
        RECT 98.260 153.325 98.430 153.825 ;
        RECT 97.400 153.035 98.090 153.205 ;
        RECT 97.400 152.445 98.090 152.615 ;
        RECT 97.060 151.825 97.230 152.325 ;
        RECT 98.260 151.825 98.430 152.325 ;
        RECT 97.400 151.535 98.090 151.705 ;
        RECT 97.400 150.945 98.090 151.115 ;
        RECT 97.060 150.325 97.230 150.825 ;
        RECT 98.260 150.325 98.430 150.825 ;
        RECT 97.400 150.035 98.090 150.205 ;
        RECT 97.400 149.445 98.090 149.615 ;
        RECT 97.060 148.825 97.230 149.325 ;
        RECT 98.260 148.825 98.430 149.325 ;
        RECT 97.400 148.535 98.090 148.705 ;
        RECT 97.400 147.945 98.090 148.115 ;
        RECT 97.060 147.325 97.230 147.825 ;
        RECT 98.260 147.325 98.430 147.825 ;
        RECT 97.400 147.035 98.090 147.205 ;
        RECT 97.400 146.445 98.090 146.615 ;
        RECT 97.060 145.825 97.230 146.325 ;
        RECT 98.260 145.825 98.430 146.325 ;
        RECT 97.400 145.535 98.090 145.705 ;
        RECT 97.400 144.945 98.090 145.115 ;
        RECT 97.060 144.325 97.230 144.825 ;
        RECT 98.260 144.325 98.430 144.825 ;
        RECT 97.400 144.035 98.090 144.205 ;
        RECT 97.400 143.445 98.090 143.615 ;
        RECT 97.060 142.825 97.230 143.325 ;
        RECT 98.260 142.825 98.430 143.325 ;
        RECT 97.400 142.535 98.090 142.705 ;
        RECT 97.400 141.945 98.090 142.115 ;
        RECT 97.060 141.325 97.230 141.825 ;
        RECT 98.260 141.325 98.430 141.825 ;
        RECT 97.400 141.035 98.090 141.205 ;
        RECT 98.725 140.495 98.895 154.605 ;
        RECT 96.595 140.325 98.895 140.495 ;
        RECT 99.775 154.505 102.425 154.675 ;
        RECT 99.775 140.645 99.945 154.505 ;
        RECT 100.580 153.945 101.620 154.115 ;
        RECT 100.195 153.325 100.365 153.825 ;
        RECT 101.835 153.325 102.005 153.825 ;
        RECT 100.580 153.035 101.620 153.205 ;
        RECT 100.580 152.445 101.620 152.615 ;
        RECT 100.195 151.825 100.365 152.325 ;
        RECT 101.835 151.825 102.005 152.325 ;
        RECT 100.580 151.535 101.620 151.705 ;
        RECT 100.580 150.945 101.620 151.115 ;
        RECT 100.195 150.325 100.365 150.825 ;
        RECT 101.835 150.325 102.005 150.825 ;
        RECT 100.580 150.035 101.620 150.205 ;
        RECT 100.580 149.445 101.620 149.615 ;
        RECT 100.195 148.825 100.365 149.325 ;
        RECT 101.835 148.825 102.005 149.325 ;
        RECT 100.580 148.535 101.620 148.705 ;
        RECT 100.580 147.945 101.620 148.115 ;
        RECT 100.195 147.325 100.365 147.825 ;
        RECT 101.835 147.325 102.005 147.825 ;
        RECT 100.580 147.035 101.620 147.205 ;
        RECT 100.580 146.445 101.620 146.615 ;
        RECT 100.195 145.825 100.365 146.325 ;
        RECT 101.835 145.825 102.005 146.325 ;
        RECT 100.580 145.535 101.620 145.705 ;
        RECT 100.580 144.945 101.620 145.115 ;
        RECT 100.195 144.325 100.365 144.825 ;
        RECT 101.835 144.325 102.005 144.825 ;
        RECT 100.580 144.035 101.620 144.205 ;
        RECT 100.580 143.445 101.620 143.615 ;
        RECT 100.195 142.825 100.365 143.325 ;
        RECT 101.835 142.825 102.005 143.325 ;
        RECT 100.580 142.535 101.620 142.705 ;
        RECT 100.580 141.945 101.620 142.115 ;
        RECT 100.195 141.325 100.365 141.825 ;
        RECT 101.835 141.325 102.005 141.825 ;
        RECT 100.580 141.035 101.620 141.205 ;
        RECT 102.255 140.645 102.425 154.505 ;
        RECT 99.775 140.475 102.425 140.645 ;
        RECT 55.745 132.745 82.915 132.915 ;
        RECT 55.745 132.435 55.915 132.745 ;
        RECT 55.550 129.355 56.050 132.435 ;
        RECT 56.685 132.280 57.185 132.450 ;
        RECT 58.065 132.280 58.565 132.450 ;
        RECT 59.445 132.280 59.945 132.450 ;
        RECT 60.825 132.280 61.325 132.450 ;
        RECT 62.205 132.280 62.705 132.450 ;
        RECT 63.585 132.280 64.085 132.450 ;
        RECT 64.965 132.280 65.465 132.450 ;
        RECT 66.345 132.280 66.845 132.450 ;
        RECT 67.725 132.280 68.225 132.450 ;
        RECT 69.105 132.280 69.605 132.450 ;
        RECT 70.485 132.280 70.985 132.450 ;
        RECT 71.865 132.280 72.365 132.450 ;
        RECT 73.245 132.280 73.745 132.450 ;
        RECT 74.625 132.280 75.125 132.450 ;
        RECT 76.005 132.280 76.505 132.450 ;
        RECT 77.385 132.280 77.885 132.450 ;
        RECT 78.765 132.280 79.265 132.450 ;
        RECT 80.145 132.280 80.645 132.450 ;
        RECT 81.525 132.280 82.025 132.450 ;
        RECT 82.745 132.435 82.915 132.745 ;
        RECT 56.455 131.420 56.625 132.110 ;
        RECT 57.245 131.420 57.415 132.110 ;
        RECT 57.835 131.420 58.005 132.110 ;
        RECT 58.625 131.420 58.795 132.110 ;
        RECT 59.215 131.420 59.385 132.110 ;
        RECT 60.005 131.420 60.175 132.110 ;
        RECT 60.595 131.420 60.765 132.110 ;
        RECT 61.385 131.420 61.555 132.110 ;
        RECT 61.975 131.420 62.145 132.110 ;
        RECT 62.765 131.420 62.935 132.110 ;
        RECT 63.355 131.420 63.525 132.110 ;
        RECT 64.145 131.420 64.315 132.110 ;
        RECT 64.735 131.420 64.905 132.110 ;
        RECT 65.525 131.420 65.695 132.110 ;
        RECT 66.115 131.420 66.285 132.110 ;
        RECT 66.905 131.420 67.075 132.110 ;
        RECT 67.495 131.420 67.665 132.110 ;
        RECT 68.285 131.420 68.455 132.110 ;
        RECT 68.875 131.420 69.045 132.110 ;
        RECT 69.665 131.420 69.835 132.110 ;
        RECT 70.255 131.420 70.425 132.110 ;
        RECT 71.045 131.420 71.215 132.110 ;
        RECT 71.635 131.420 71.805 132.110 ;
        RECT 72.425 131.420 72.595 132.110 ;
        RECT 73.015 131.420 73.185 132.110 ;
        RECT 73.805 131.420 73.975 132.110 ;
        RECT 74.395 131.420 74.565 132.110 ;
        RECT 75.185 131.420 75.355 132.110 ;
        RECT 75.775 131.420 75.945 132.110 ;
        RECT 76.565 131.420 76.735 132.110 ;
        RECT 77.155 131.420 77.325 132.110 ;
        RECT 77.945 131.420 78.115 132.110 ;
        RECT 78.535 131.420 78.705 132.110 ;
        RECT 79.325 131.420 79.495 132.110 ;
        RECT 79.915 131.420 80.085 132.110 ;
        RECT 80.705 131.420 80.875 132.110 ;
        RECT 81.295 131.420 81.465 132.110 ;
        RECT 82.085 131.420 82.255 132.110 ;
        RECT 56.685 131.080 57.185 131.250 ;
        RECT 58.065 131.080 58.565 131.250 ;
        RECT 59.445 131.080 59.945 131.250 ;
        RECT 60.825 131.080 61.325 131.250 ;
        RECT 62.205 131.080 62.705 131.250 ;
        RECT 63.585 131.080 64.085 131.250 ;
        RECT 64.965 131.080 65.465 131.250 ;
        RECT 66.345 131.080 66.845 131.250 ;
        RECT 67.725 131.080 68.225 131.250 ;
        RECT 69.105 131.080 69.605 131.250 ;
        RECT 70.485 131.080 70.985 131.250 ;
        RECT 71.865 131.080 72.365 131.250 ;
        RECT 73.245 131.080 73.745 131.250 ;
        RECT 74.625 131.080 75.125 131.250 ;
        RECT 76.005 131.080 76.505 131.250 ;
        RECT 77.385 131.080 77.885 131.250 ;
        RECT 78.765 131.080 79.265 131.250 ;
        RECT 80.145 131.080 80.645 131.250 ;
        RECT 81.525 131.080 82.025 131.250 ;
        RECT 56.685 130.540 57.185 130.710 ;
        RECT 58.065 130.540 58.565 130.710 ;
        RECT 59.445 130.540 59.945 130.710 ;
        RECT 60.825 130.540 61.325 130.710 ;
        RECT 62.205 130.540 62.705 130.710 ;
        RECT 63.585 130.540 64.085 130.710 ;
        RECT 64.965 130.540 65.465 130.710 ;
        RECT 66.345 130.540 66.845 130.710 ;
        RECT 67.725 130.540 68.225 130.710 ;
        RECT 69.105 130.540 69.605 130.710 ;
        RECT 70.485 130.540 70.985 130.710 ;
        RECT 71.865 130.540 72.365 130.710 ;
        RECT 73.245 130.540 73.745 130.710 ;
        RECT 74.625 130.540 75.125 130.710 ;
        RECT 76.005 130.540 76.505 130.710 ;
        RECT 77.385 130.540 77.885 130.710 ;
        RECT 78.765 130.540 79.265 130.710 ;
        RECT 80.145 130.540 80.645 130.710 ;
        RECT 81.525 130.540 82.025 130.710 ;
        RECT 56.455 129.680 56.625 130.370 ;
        RECT 57.245 129.680 57.415 130.370 ;
        RECT 57.835 129.680 58.005 130.370 ;
        RECT 58.625 129.680 58.795 130.370 ;
        RECT 59.215 129.680 59.385 130.370 ;
        RECT 60.005 129.680 60.175 130.370 ;
        RECT 60.595 129.680 60.765 130.370 ;
        RECT 61.385 129.680 61.555 130.370 ;
        RECT 61.975 129.680 62.145 130.370 ;
        RECT 62.765 129.680 62.935 130.370 ;
        RECT 63.355 129.680 63.525 130.370 ;
        RECT 64.145 129.680 64.315 130.370 ;
        RECT 64.735 129.680 64.905 130.370 ;
        RECT 65.525 129.680 65.695 130.370 ;
        RECT 66.115 129.680 66.285 130.370 ;
        RECT 66.905 129.680 67.075 130.370 ;
        RECT 67.495 129.680 67.665 130.370 ;
        RECT 68.285 129.680 68.455 130.370 ;
        RECT 68.875 129.680 69.045 130.370 ;
        RECT 69.665 129.680 69.835 130.370 ;
        RECT 70.255 129.680 70.425 130.370 ;
        RECT 71.045 129.680 71.215 130.370 ;
        RECT 71.635 129.680 71.805 130.370 ;
        RECT 72.425 129.680 72.595 130.370 ;
        RECT 73.015 129.680 73.185 130.370 ;
        RECT 73.805 129.680 73.975 130.370 ;
        RECT 74.395 129.680 74.565 130.370 ;
        RECT 75.185 129.680 75.355 130.370 ;
        RECT 75.775 129.680 75.945 130.370 ;
        RECT 76.565 129.680 76.735 130.370 ;
        RECT 77.155 129.680 77.325 130.370 ;
        RECT 77.945 129.680 78.115 130.370 ;
        RECT 78.535 129.680 78.705 130.370 ;
        RECT 79.325 129.680 79.495 130.370 ;
        RECT 79.915 129.680 80.085 130.370 ;
        RECT 80.705 129.680 80.875 130.370 ;
        RECT 81.295 129.680 81.465 130.370 ;
        RECT 82.085 129.680 82.255 130.370 ;
        RECT 55.745 129.045 55.915 129.355 ;
        RECT 56.685 129.340 57.185 129.510 ;
        RECT 58.065 129.340 58.565 129.510 ;
        RECT 59.445 129.340 59.945 129.510 ;
        RECT 60.825 129.340 61.325 129.510 ;
        RECT 62.205 129.340 62.705 129.510 ;
        RECT 63.585 129.340 64.085 129.510 ;
        RECT 64.965 129.340 65.465 129.510 ;
        RECT 66.345 129.340 66.845 129.510 ;
        RECT 67.725 129.340 68.225 129.510 ;
        RECT 69.105 129.340 69.605 129.510 ;
        RECT 70.485 129.340 70.985 129.510 ;
        RECT 71.865 129.340 72.365 129.510 ;
        RECT 73.245 129.340 73.745 129.510 ;
        RECT 74.625 129.340 75.125 129.510 ;
        RECT 76.005 129.340 76.505 129.510 ;
        RECT 77.385 129.340 77.885 129.510 ;
        RECT 78.765 129.340 79.265 129.510 ;
        RECT 80.145 129.340 80.645 129.510 ;
        RECT 81.525 129.340 82.025 129.510 ;
        RECT 82.660 129.355 83.160 132.435 ;
        RECT 82.745 129.045 82.915 129.355 ;
        RECT 55.745 128.875 82.915 129.045 ;
        RECT 55.895 127.825 82.815 127.995 ;
        RECT 55.895 127.515 56.065 127.825 ;
        RECT 55.550 123.335 56.065 127.515 ;
        RECT 56.685 127.405 57.185 127.575 ;
        RECT 58.065 127.405 58.565 127.575 ;
        RECT 59.445 127.405 59.945 127.575 ;
        RECT 60.825 127.405 61.325 127.575 ;
        RECT 62.205 127.405 62.705 127.575 ;
        RECT 63.585 127.405 64.085 127.575 ;
        RECT 64.965 127.405 65.465 127.575 ;
        RECT 66.345 127.405 66.845 127.575 ;
        RECT 67.725 127.405 68.225 127.575 ;
        RECT 69.105 127.405 69.605 127.575 ;
        RECT 70.485 127.405 70.985 127.575 ;
        RECT 71.865 127.405 72.365 127.575 ;
        RECT 73.245 127.405 73.745 127.575 ;
        RECT 74.625 127.405 75.125 127.575 ;
        RECT 76.005 127.405 76.505 127.575 ;
        RECT 77.385 127.405 77.885 127.575 ;
        RECT 78.765 127.405 79.265 127.575 ;
        RECT 80.145 127.405 80.645 127.575 ;
        RECT 81.525 127.405 82.025 127.575 ;
        RECT 82.645 127.515 82.815 127.825 ;
        RECT 56.455 126.150 56.625 127.190 ;
        RECT 57.245 126.150 57.415 127.190 ;
        RECT 57.835 126.150 58.005 127.190 ;
        RECT 58.625 126.150 58.795 127.190 ;
        RECT 59.215 126.150 59.385 127.190 ;
        RECT 60.005 126.150 60.175 127.190 ;
        RECT 60.595 126.150 60.765 127.190 ;
        RECT 61.385 126.150 61.555 127.190 ;
        RECT 61.975 126.150 62.145 127.190 ;
        RECT 62.765 126.150 62.935 127.190 ;
        RECT 63.355 126.150 63.525 127.190 ;
        RECT 64.145 126.150 64.315 127.190 ;
        RECT 64.735 126.150 64.905 127.190 ;
        RECT 65.525 126.150 65.695 127.190 ;
        RECT 66.115 126.150 66.285 127.190 ;
        RECT 66.905 126.150 67.075 127.190 ;
        RECT 67.495 126.150 67.665 127.190 ;
        RECT 68.285 126.150 68.455 127.190 ;
        RECT 68.875 126.150 69.045 127.190 ;
        RECT 69.665 126.150 69.835 127.190 ;
        RECT 70.255 126.150 70.425 127.190 ;
        RECT 71.045 126.150 71.215 127.190 ;
        RECT 71.635 126.150 71.805 127.190 ;
        RECT 72.425 126.150 72.595 127.190 ;
        RECT 73.015 126.150 73.185 127.190 ;
        RECT 73.805 126.150 73.975 127.190 ;
        RECT 74.395 126.150 74.565 127.190 ;
        RECT 75.185 126.150 75.355 127.190 ;
        RECT 75.775 126.150 75.945 127.190 ;
        RECT 76.565 126.150 76.735 127.190 ;
        RECT 77.155 126.150 77.325 127.190 ;
        RECT 77.945 126.150 78.115 127.190 ;
        RECT 78.535 126.150 78.705 127.190 ;
        RECT 79.325 126.150 79.495 127.190 ;
        RECT 79.915 126.150 80.085 127.190 ;
        RECT 80.705 126.150 80.875 127.190 ;
        RECT 81.295 126.150 81.465 127.190 ;
        RECT 82.085 126.150 82.255 127.190 ;
        RECT 56.685 125.765 57.185 125.935 ;
        RECT 58.065 125.765 58.565 125.935 ;
        RECT 59.445 125.765 59.945 125.935 ;
        RECT 60.825 125.765 61.325 125.935 ;
        RECT 62.205 125.765 62.705 125.935 ;
        RECT 63.585 125.765 64.085 125.935 ;
        RECT 64.965 125.765 65.465 125.935 ;
        RECT 66.345 125.765 66.845 125.935 ;
        RECT 67.725 125.765 68.225 125.935 ;
        RECT 69.105 125.765 69.605 125.935 ;
        RECT 70.485 125.765 70.985 125.935 ;
        RECT 71.865 125.765 72.365 125.935 ;
        RECT 73.245 125.765 73.745 125.935 ;
        RECT 74.625 125.765 75.125 125.935 ;
        RECT 76.005 125.765 76.505 125.935 ;
        RECT 77.385 125.765 77.885 125.935 ;
        RECT 78.765 125.765 79.265 125.935 ;
        RECT 80.145 125.765 80.645 125.935 ;
        RECT 81.525 125.765 82.025 125.935 ;
        RECT 56.685 125.225 57.185 125.395 ;
        RECT 58.065 125.225 58.565 125.395 ;
        RECT 59.445 125.225 59.945 125.395 ;
        RECT 60.825 125.225 61.325 125.395 ;
        RECT 62.205 125.225 62.705 125.395 ;
        RECT 63.585 125.225 64.085 125.395 ;
        RECT 64.965 125.225 65.465 125.395 ;
        RECT 66.345 125.225 66.845 125.395 ;
        RECT 67.725 125.225 68.225 125.395 ;
        RECT 69.105 125.225 69.605 125.395 ;
        RECT 70.485 125.225 70.985 125.395 ;
        RECT 71.865 125.225 72.365 125.395 ;
        RECT 73.245 125.225 73.745 125.395 ;
        RECT 74.625 125.225 75.125 125.395 ;
        RECT 76.005 125.225 76.505 125.395 ;
        RECT 77.385 125.225 77.885 125.395 ;
        RECT 78.765 125.225 79.265 125.395 ;
        RECT 80.145 125.225 80.645 125.395 ;
        RECT 81.525 125.225 82.025 125.395 ;
        RECT 56.455 123.970 56.625 125.010 ;
        RECT 57.245 123.970 57.415 125.010 ;
        RECT 57.835 123.970 58.005 125.010 ;
        RECT 58.625 123.970 58.795 125.010 ;
        RECT 59.215 123.970 59.385 125.010 ;
        RECT 60.005 123.970 60.175 125.010 ;
        RECT 60.595 123.970 60.765 125.010 ;
        RECT 61.385 123.970 61.555 125.010 ;
        RECT 61.975 123.970 62.145 125.010 ;
        RECT 62.765 123.970 62.935 125.010 ;
        RECT 63.355 123.970 63.525 125.010 ;
        RECT 64.145 123.970 64.315 125.010 ;
        RECT 64.735 123.970 64.905 125.010 ;
        RECT 65.525 123.970 65.695 125.010 ;
        RECT 66.115 123.970 66.285 125.010 ;
        RECT 66.905 123.970 67.075 125.010 ;
        RECT 67.495 123.970 67.665 125.010 ;
        RECT 68.285 123.970 68.455 125.010 ;
        RECT 68.875 123.970 69.045 125.010 ;
        RECT 69.665 123.970 69.835 125.010 ;
        RECT 70.255 123.970 70.425 125.010 ;
        RECT 71.045 123.970 71.215 125.010 ;
        RECT 71.635 123.970 71.805 125.010 ;
        RECT 72.425 123.970 72.595 125.010 ;
        RECT 73.015 123.970 73.185 125.010 ;
        RECT 73.805 123.970 73.975 125.010 ;
        RECT 74.395 123.970 74.565 125.010 ;
        RECT 75.185 123.970 75.355 125.010 ;
        RECT 75.775 123.970 75.945 125.010 ;
        RECT 76.565 123.970 76.735 125.010 ;
        RECT 77.155 123.970 77.325 125.010 ;
        RECT 77.945 123.970 78.115 125.010 ;
        RECT 78.535 123.970 78.705 125.010 ;
        RECT 79.325 123.970 79.495 125.010 ;
        RECT 79.915 123.970 80.085 125.010 ;
        RECT 80.705 123.970 80.875 125.010 ;
        RECT 81.295 123.970 81.465 125.010 ;
        RECT 82.085 123.970 82.255 125.010 ;
        RECT 56.685 123.585 57.185 123.755 ;
        RECT 58.065 123.585 58.565 123.755 ;
        RECT 59.445 123.585 59.945 123.755 ;
        RECT 60.825 123.585 61.325 123.755 ;
        RECT 62.205 123.585 62.705 123.755 ;
        RECT 63.585 123.585 64.085 123.755 ;
        RECT 64.965 123.585 65.465 123.755 ;
        RECT 66.345 123.585 66.845 123.755 ;
        RECT 67.725 123.585 68.225 123.755 ;
        RECT 69.105 123.585 69.605 123.755 ;
        RECT 70.485 123.585 70.985 123.755 ;
        RECT 71.865 123.585 72.365 123.755 ;
        RECT 73.245 123.585 73.745 123.755 ;
        RECT 74.625 123.585 75.125 123.755 ;
        RECT 76.005 123.585 76.505 123.755 ;
        RECT 77.385 123.585 77.885 123.755 ;
        RECT 78.765 123.585 79.265 123.755 ;
        RECT 80.145 123.585 80.645 123.755 ;
        RECT 81.525 123.585 82.025 123.755 ;
        RECT 82.645 123.335 83.160 127.515 ;
        RECT 55.550 123.190 83.160 123.335 ;
        RECT 55.895 123.165 82.815 123.190 ;
        RECT 55.190 121.660 83.520 121.830 ;
        RECT 55.190 121.350 55.360 121.660 ;
        RECT 54.800 107.980 55.360 121.350 ;
        RECT 83.350 121.350 83.520 121.660 ;
        RECT 55.900 118.960 56.250 121.120 ;
        RECT 56.730 118.960 57.080 121.120 ;
        RECT 57.560 118.960 57.910 121.120 ;
        RECT 58.390 118.960 58.740 121.120 ;
        RECT 59.220 118.960 59.570 121.120 ;
        RECT 60.050 118.960 60.400 121.120 ;
        RECT 60.880 118.960 61.230 121.120 ;
        RECT 61.710 118.960 62.060 121.120 ;
        RECT 62.540 118.960 62.890 121.120 ;
        RECT 63.370 118.960 63.720 121.120 ;
        RECT 64.200 118.960 64.550 121.120 ;
        RECT 65.030 118.960 65.380 121.120 ;
        RECT 65.860 118.960 66.210 121.120 ;
        RECT 66.690 118.960 67.040 121.120 ;
        RECT 67.520 118.960 67.870 121.120 ;
        RECT 68.350 118.960 68.700 121.120 ;
        RECT 69.180 118.960 69.530 121.120 ;
        RECT 70.010 118.960 70.360 121.120 ;
        RECT 70.840 118.960 71.190 121.120 ;
        RECT 71.670 118.960 72.020 121.120 ;
        RECT 72.500 118.960 72.850 121.120 ;
        RECT 73.330 118.960 73.680 121.120 ;
        RECT 74.160 118.960 74.510 121.120 ;
        RECT 74.990 118.960 75.340 121.120 ;
        RECT 75.820 118.960 76.170 121.120 ;
        RECT 76.650 118.960 77.000 121.120 ;
        RECT 77.480 118.960 77.830 121.120 ;
        RECT 78.310 118.960 78.660 121.120 ;
        RECT 79.140 118.960 79.490 121.120 ;
        RECT 79.970 118.960 80.320 121.120 ;
        RECT 80.800 118.960 81.150 121.120 ;
        RECT 81.630 118.960 81.980 121.120 ;
        RECT 82.460 118.960 82.810 121.120 ;
        RECT 55.900 108.210 56.250 110.370 ;
        RECT 56.730 108.210 57.080 110.370 ;
        RECT 57.560 108.210 57.910 110.370 ;
        RECT 58.390 108.210 58.740 110.370 ;
        RECT 59.220 108.210 59.570 110.370 ;
        RECT 60.050 108.210 60.400 110.370 ;
        RECT 60.880 108.210 61.230 110.370 ;
        RECT 61.710 108.210 62.060 110.370 ;
        RECT 62.540 108.210 62.890 110.370 ;
        RECT 63.370 108.210 63.720 110.370 ;
        RECT 64.200 108.210 64.550 110.370 ;
        RECT 65.030 108.210 65.380 110.370 ;
        RECT 65.860 108.210 66.210 110.370 ;
        RECT 66.690 108.210 67.040 110.370 ;
        RECT 67.520 108.210 67.870 110.370 ;
        RECT 68.350 108.210 68.700 110.370 ;
        RECT 69.180 108.210 69.530 110.370 ;
        RECT 70.010 108.210 70.360 110.370 ;
        RECT 70.840 108.210 71.190 110.370 ;
        RECT 71.670 108.210 72.020 110.370 ;
        RECT 72.500 108.210 72.850 110.370 ;
        RECT 73.330 108.210 73.680 110.370 ;
        RECT 74.160 108.210 74.510 110.370 ;
        RECT 74.990 108.210 75.340 110.370 ;
        RECT 75.820 108.210 76.170 110.370 ;
        RECT 76.650 108.210 77.000 110.370 ;
        RECT 77.480 108.210 77.830 110.370 ;
        RECT 78.310 108.210 78.660 110.370 ;
        RECT 79.140 108.210 79.490 110.370 ;
        RECT 79.970 108.210 80.320 110.370 ;
        RECT 80.800 108.210 81.150 110.370 ;
        RECT 81.630 108.210 81.980 110.370 ;
        RECT 82.460 108.210 82.810 110.370 ;
        RECT 55.190 107.670 55.360 107.980 ;
        RECT 83.350 107.980 83.910 121.350 ;
        RECT 83.350 107.670 83.520 107.980 ;
        RECT 55.190 107.500 83.520 107.670 ;
        RECT 55.895 106.140 82.815 106.165 ;
        RECT 55.550 105.995 83.160 106.140 ;
        RECT 55.550 101.815 56.065 105.995 ;
        RECT 56.685 105.575 57.185 105.745 ;
        RECT 58.065 105.575 58.565 105.745 ;
        RECT 59.445 105.575 59.945 105.745 ;
        RECT 60.825 105.575 61.325 105.745 ;
        RECT 62.205 105.575 62.705 105.745 ;
        RECT 63.585 105.575 64.085 105.745 ;
        RECT 64.965 105.575 65.465 105.745 ;
        RECT 66.345 105.575 66.845 105.745 ;
        RECT 67.725 105.575 68.225 105.745 ;
        RECT 69.105 105.575 69.605 105.745 ;
        RECT 70.485 105.575 70.985 105.745 ;
        RECT 71.865 105.575 72.365 105.745 ;
        RECT 73.245 105.575 73.745 105.745 ;
        RECT 74.625 105.575 75.125 105.745 ;
        RECT 76.005 105.575 76.505 105.745 ;
        RECT 77.385 105.575 77.885 105.745 ;
        RECT 78.765 105.575 79.265 105.745 ;
        RECT 80.145 105.575 80.645 105.745 ;
        RECT 81.525 105.575 82.025 105.745 ;
        RECT 56.455 104.320 56.625 105.360 ;
        RECT 57.245 104.320 57.415 105.360 ;
        RECT 57.835 104.320 58.005 105.360 ;
        RECT 58.625 104.320 58.795 105.360 ;
        RECT 59.215 104.320 59.385 105.360 ;
        RECT 60.005 104.320 60.175 105.360 ;
        RECT 60.595 104.320 60.765 105.360 ;
        RECT 61.385 104.320 61.555 105.360 ;
        RECT 61.975 104.320 62.145 105.360 ;
        RECT 62.765 104.320 62.935 105.360 ;
        RECT 63.355 104.320 63.525 105.360 ;
        RECT 64.145 104.320 64.315 105.360 ;
        RECT 64.735 104.320 64.905 105.360 ;
        RECT 65.525 104.320 65.695 105.360 ;
        RECT 66.115 104.320 66.285 105.360 ;
        RECT 66.905 104.320 67.075 105.360 ;
        RECT 67.495 104.320 67.665 105.360 ;
        RECT 68.285 104.320 68.455 105.360 ;
        RECT 68.875 104.320 69.045 105.360 ;
        RECT 69.665 104.320 69.835 105.360 ;
        RECT 70.255 104.320 70.425 105.360 ;
        RECT 71.045 104.320 71.215 105.360 ;
        RECT 71.635 104.320 71.805 105.360 ;
        RECT 72.425 104.320 72.595 105.360 ;
        RECT 73.015 104.320 73.185 105.360 ;
        RECT 73.805 104.320 73.975 105.360 ;
        RECT 74.395 104.320 74.565 105.360 ;
        RECT 75.185 104.320 75.355 105.360 ;
        RECT 75.775 104.320 75.945 105.360 ;
        RECT 76.565 104.320 76.735 105.360 ;
        RECT 77.155 104.320 77.325 105.360 ;
        RECT 77.945 104.320 78.115 105.360 ;
        RECT 78.535 104.320 78.705 105.360 ;
        RECT 79.325 104.320 79.495 105.360 ;
        RECT 79.915 104.320 80.085 105.360 ;
        RECT 80.705 104.320 80.875 105.360 ;
        RECT 81.295 104.320 81.465 105.360 ;
        RECT 82.085 104.320 82.255 105.360 ;
        RECT 56.685 103.935 57.185 104.105 ;
        RECT 58.065 103.935 58.565 104.105 ;
        RECT 59.445 103.935 59.945 104.105 ;
        RECT 60.825 103.935 61.325 104.105 ;
        RECT 62.205 103.935 62.705 104.105 ;
        RECT 63.585 103.935 64.085 104.105 ;
        RECT 64.965 103.935 65.465 104.105 ;
        RECT 66.345 103.935 66.845 104.105 ;
        RECT 67.725 103.935 68.225 104.105 ;
        RECT 69.105 103.935 69.605 104.105 ;
        RECT 70.485 103.935 70.985 104.105 ;
        RECT 71.865 103.935 72.365 104.105 ;
        RECT 73.245 103.935 73.745 104.105 ;
        RECT 74.625 103.935 75.125 104.105 ;
        RECT 76.005 103.935 76.505 104.105 ;
        RECT 77.385 103.935 77.885 104.105 ;
        RECT 78.765 103.935 79.265 104.105 ;
        RECT 80.145 103.935 80.645 104.105 ;
        RECT 81.525 103.935 82.025 104.105 ;
        RECT 56.685 103.395 57.185 103.565 ;
        RECT 58.065 103.395 58.565 103.565 ;
        RECT 59.445 103.395 59.945 103.565 ;
        RECT 60.825 103.395 61.325 103.565 ;
        RECT 62.205 103.395 62.705 103.565 ;
        RECT 63.585 103.395 64.085 103.565 ;
        RECT 64.965 103.395 65.465 103.565 ;
        RECT 66.345 103.395 66.845 103.565 ;
        RECT 67.725 103.395 68.225 103.565 ;
        RECT 69.105 103.395 69.605 103.565 ;
        RECT 70.485 103.395 70.985 103.565 ;
        RECT 71.865 103.395 72.365 103.565 ;
        RECT 73.245 103.395 73.745 103.565 ;
        RECT 74.625 103.395 75.125 103.565 ;
        RECT 76.005 103.395 76.505 103.565 ;
        RECT 77.385 103.395 77.885 103.565 ;
        RECT 78.765 103.395 79.265 103.565 ;
        RECT 80.145 103.395 80.645 103.565 ;
        RECT 81.525 103.395 82.025 103.565 ;
        RECT 56.455 102.140 56.625 103.180 ;
        RECT 57.245 102.140 57.415 103.180 ;
        RECT 57.835 102.140 58.005 103.180 ;
        RECT 58.625 102.140 58.795 103.180 ;
        RECT 59.215 102.140 59.385 103.180 ;
        RECT 60.005 102.140 60.175 103.180 ;
        RECT 60.595 102.140 60.765 103.180 ;
        RECT 61.385 102.140 61.555 103.180 ;
        RECT 61.975 102.140 62.145 103.180 ;
        RECT 62.765 102.140 62.935 103.180 ;
        RECT 63.355 102.140 63.525 103.180 ;
        RECT 64.145 102.140 64.315 103.180 ;
        RECT 64.735 102.140 64.905 103.180 ;
        RECT 65.525 102.140 65.695 103.180 ;
        RECT 66.115 102.140 66.285 103.180 ;
        RECT 66.905 102.140 67.075 103.180 ;
        RECT 67.495 102.140 67.665 103.180 ;
        RECT 68.285 102.140 68.455 103.180 ;
        RECT 68.875 102.140 69.045 103.180 ;
        RECT 69.665 102.140 69.835 103.180 ;
        RECT 70.255 102.140 70.425 103.180 ;
        RECT 71.045 102.140 71.215 103.180 ;
        RECT 71.635 102.140 71.805 103.180 ;
        RECT 72.425 102.140 72.595 103.180 ;
        RECT 73.015 102.140 73.185 103.180 ;
        RECT 73.805 102.140 73.975 103.180 ;
        RECT 74.395 102.140 74.565 103.180 ;
        RECT 75.185 102.140 75.355 103.180 ;
        RECT 75.775 102.140 75.945 103.180 ;
        RECT 76.565 102.140 76.735 103.180 ;
        RECT 77.155 102.140 77.325 103.180 ;
        RECT 77.945 102.140 78.115 103.180 ;
        RECT 78.535 102.140 78.705 103.180 ;
        RECT 79.325 102.140 79.495 103.180 ;
        RECT 79.915 102.140 80.085 103.180 ;
        RECT 80.705 102.140 80.875 103.180 ;
        RECT 81.295 102.140 81.465 103.180 ;
        RECT 82.085 102.140 82.255 103.180 ;
        RECT 55.895 101.505 56.065 101.815 ;
        RECT 56.685 101.755 57.185 101.925 ;
        RECT 58.065 101.755 58.565 101.925 ;
        RECT 59.445 101.755 59.945 101.925 ;
        RECT 60.825 101.755 61.325 101.925 ;
        RECT 62.205 101.755 62.705 101.925 ;
        RECT 63.585 101.755 64.085 101.925 ;
        RECT 64.965 101.755 65.465 101.925 ;
        RECT 66.345 101.755 66.845 101.925 ;
        RECT 67.725 101.755 68.225 101.925 ;
        RECT 69.105 101.755 69.605 101.925 ;
        RECT 70.485 101.755 70.985 101.925 ;
        RECT 71.865 101.755 72.365 101.925 ;
        RECT 73.245 101.755 73.745 101.925 ;
        RECT 74.625 101.755 75.125 101.925 ;
        RECT 76.005 101.755 76.505 101.925 ;
        RECT 77.385 101.755 77.885 101.925 ;
        RECT 78.765 101.755 79.265 101.925 ;
        RECT 80.145 101.755 80.645 101.925 ;
        RECT 81.525 101.755 82.025 101.925 ;
        RECT 82.645 101.815 83.160 105.995 ;
        RECT 82.645 101.505 82.815 101.815 ;
        RECT 55.895 101.335 82.815 101.505 ;
        RECT 55.795 100.285 82.965 100.455 ;
        RECT 55.795 99.975 55.965 100.285 ;
        RECT 55.550 96.895 56.050 99.975 ;
        RECT 56.685 99.820 57.185 99.990 ;
        RECT 58.065 99.820 58.565 99.990 ;
        RECT 59.445 99.820 59.945 99.990 ;
        RECT 60.825 99.820 61.325 99.990 ;
        RECT 62.205 99.820 62.705 99.990 ;
        RECT 63.585 99.820 64.085 99.990 ;
        RECT 64.965 99.820 65.465 99.990 ;
        RECT 66.345 99.820 66.845 99.990 ;
        RECT 67.725 99.820 68.225 99.990 ;
        RECT 69.105 99.820 69.605 99.990 ;
        RECT 70.485 99.820 70.985 99.990 ;
        RECT 71.865 99.820 72.365 99.990 ;
        RECT 73.245 99.820 73.745 99.990 ;
        RECT 74.625 99.820 75.125 99.990 ;
        RECT 76.005 99.820 76.505 99.990 ;
        RECT 77.385 99.820 77.885 99.990 ;
        RECT 78.765 99.820 79.265 99.990 ;
        RECT 80.145 99.820 80.645 99.990 ;
        RECT 81.525 99.820 82.025 99.990 ;
        RECT 82.795 99.975 82.965 100.285 ;
        RECT 56.455 98.960 56.625 99.650 ;
        RECT 57.245 98.960 57.415 99.650 ;
        RECT 57.835 98.960 58.005 99.650 ;
        RECT 58.625 98.960 58.795 99.650 ;
        RECT 59.215 98.960 59.385 99.650 ;
        RECT 60.005 98.960 60.175 99.650 ;
        RECT 60.595 98.960 60.765 99.650 ;
        RECT 61.385 98.960 61.555 99.650 ;
        RECT 61.975 98.960 62.145 99.650 ;
        RECT 62.765 98.960 62.935 99.650 ;
        RECT 63.355 98.960 63.525 99.650 ;
        RECT 64.145 98.960 64.315 99.650 ;
        RECT 64.735 98.960 64.905 99.650 ;
        RECT 65.525 98.960 65.695 99.650 ;
        RECT 66.115 98.960 66.285 99.650 ;
        RECT 66.905 98.960 67.075 99.650 ;
        RECT 67.495 98.960 67.665 99.650 ;
        RECT 68.285 98.960 68.455 99.650 ;
        RECT 68.875 98.960 69.045 99.650 ;
        RECT 69.665 98.960 69.835 99.650 ;
        RECT 70.255 98.960 70.425 99.650 ;
        RECT 71.045 98.960 71.215 99.650 ;
        RECT 71.635 98.960 71.805 99.650 ;
        RECT 72.425 98.960 72.595 99.650 ;
        RECT 73.015 98.960 73.185 99.650 ;
        RECT 73.805 98.960 73.975 99.650 ;
        RECT 74.395 98.960 74.565 99.650 ;
        RECT 75.185 98.960 75.355 99.650 ;
        RECT 75.775 98.960 75.945 99.650 ;
        RECT 76.565 98.960 76.735 99.650 ;
        RECT 77.155 98.960 77.325 99.650 ;
        RECT 77.945 98.960 78.115 99.650 ;
        RECT 78.535 98.960 78.705 99.650 ;
        RECT 79.325 98.960 79.495 99.650 ;
        RECT 79.915 98.960 80.085 99.650 ;
        RECT 80.705 98.960 80.875 99.650 ;
        RECT 81.295 98.960 81.465 99.650 ;
        RECT 82.085 98.960 82.255 99.650 ;
        RECT 56.685 98.620 57.185 98.790 ;
        RECT 58.065 98.620 58.565 98.790 ;
        RECT 59.445 98.620 59.945 98.790 ;
        RECT 60.825 98.620 61.325 98.790 ;
        RECT 62.205 98.620 62.705 98.790 ;
        RECT 63.585 98.620 64.085 98.790 ;
        RECT 64.965 98.620 65.465 98.790 ;
        RECT 66.345 98.620 66.845 98.790 ;
        RECT 67.725 98.620 68.225 98.790 ;
        RECT 69.105 98.620 69.605 98.790 ;
        RECT 70.485 98.620 70.985 98.790 ;
        RECT 71.865 98.620 72.365 98.790 ;
        RECT 73.245 98.620 73.745 98.790 ;
        RECT 74.625 98.620 75.125 98.790 ;
        RECT 76.005 98.620 76.505 98.790 ;
        RECT 77.385 98.620 77.885 98.790 ;
        RECT 78.765 98.620 79.265 98.790 ;
        RECT 80.145 98.620 80.645 98.790 ;
        RECT 81.525 98.620 82.025 98.790 ;
        RECT 56.685 98.080 57.185 98.250 ;
        RECT 58.065 98.080 58.565 98.250 ;
        RECT 59.445 98.080 59.945 98.250 ;
        RECT 60.825 98.080 61.325 98.250 ;
        RECT 62.205 98.080 62.705 98.250 ;
        RECT 63.585 98.080 64.085 98.250 ;
        RECT 64.965 98.080 65.465 98.250 ;
        RECT 66.345 98.080 66.845 98.250 ;
        RECT 67.725 98.080 68.225 98.250 ;
        RECT 69.105 98.080 69.605 98.250 ;
        RECT 70.485 98.080 70.985 98.250 ;
        RECT 71.865 98.080 72.365 98.250 ;
        RECT 73.245 98.080 73.745 98.250 ;
        RECT 74.625 98.080 75.125 98.250 ;
        RECT 76.005 98.080 76.505 98.250 ;
        RECT 77.385 98.080 77.885 98.250 ;
        RECT 78.765 98.080 79.265 98.250 ;
        RECT 80.145 98.080 80.645 98.250 ;
        RECT 81.525 98.080 82.025 98.250 ;
        RECT 56.455 97.220 56.625 97.910 ;
        RECT 57.245 97.220 57.415 97.910 ;
        RECT 57.835 97.220 58.005 97.910 ;
        RECT 58.625 97.220 58.795 97.910 ;
        RECT 59.215 97.220 59.385 97.910 ;
        RECT 60.005 97.220 60.175 97.910 ;
        RECT 60.595 97.220 60.765 97.910 ;
        RECT 61.385 97.220 61.555 97.910 ;
        RECT 61.975 97.220 62.145 97.910 ;
        RECT 62.765 97.220 62.935 97.910 ;
        RECT 63.355 97.220 63.525 97.910 ;
        RECT 64.145 97.220 64.315 97.910 ;
        RECT 64.735 97.220 64.905 97.910 ;
        RECT 65.525 97.220 65.695 97.910 ;
        RECT 66.115 97.220 66.285 97.910 ;
        RECT 66.905 97.220 67.075 97.910 ;
        RECT 67.495 97.220 67.665 97.910 ;
        RECT 68.285 97.220 68.455 97.910 ;
        RECT 68.875 97.220 69.045 97.910 ;
        RECT 69.665 97.220 69.835 97.910 ;
        RECT 70.255 97.220 70.425 97.910 ;
        RECT 71.045 97.220 71.215 97.910 ;
        RECT 71.635 97.220 71.805 97.910 ;
        RECT 72.425 97.220 72.595 97.910 ;
        RECT 73.015 97.220 73.185 97.910 ;
        RECT 73.805 97.220 73.975 97.910 ;
        RECT 74.395 97.220 74.565 97.910 ;
        RECT 75.185 97.220 75.355 97.910 ;
        RECT 75.775 97.220 75.945 97.910 ;
        RECT 76.565 97.220 76.735 97.910 ;
        RECT 77.155 97.220 77.325 97.910 ;
        RECT 77.945 97.220 78.115 97.910 ;
        RECT 78.535 97.220 78.705 97.910 ;
        RECT 79.325 97.220 79.495 97.910 ;
        RECT 79.915 97.220 80.085 97.910 ;
        RECT 80.705 97.220 80.875 97.910 ;
        RECT 81.295 97.220 81.465 97.910 ;
        RECT 82.085 97.220 82.255 97.910 ;
        RECT 55.795 96.585 55.965 96.895 ;
        RECT 56.685 96.880 57.185 97.050 ;
        RECT 58.065 96.880 58.565 97.050 ;
        RECT 59.445 96.880 59.945 97.050 ;
        RECT 60.825 96.880 61.325 97.050 ;
        RECT 62.205 96.880 62.705 97.050 ;
        RECT 63.585 96.880 64.085 97.050 ;
        RECT 64.965 96.880 65.465 97.050 ;
        RECT 66.345 96.880 66.845 97.050 ;
        RECT 67.725 96.880 68.225 97.050 ;
        RECT 69.105 96.880 69.605 97.050 ;
        RECT 70.485 96.880 70.985 97.050 ;
        RECT 71.865 96.880 72.365 97.050 ;
        RECT 73.245 96.880 73.745 97.050 ;
        RECT 74.625 96.880 75.125 97.050 ;
        RECT 76.005 96.880 76.505 97.050 ;
        RECT 77.385 96.880 77.885 97.050 ;
        RECT 78.765 96.880 79.265 97.050 ;
        RECT 80.145 96.880 80.645 97.050 ;
        RECT 81.525 96.880 82.025 97.050 ;
        RECT 82.660 96.895 83.160 99.975 ;
        RECT 82.795 96.585 82.965 96.895 ;
        RECT 55.795 96.415 82.965 96.585 ;
        RECT 30.715 91.515 107.915 91.685 ;
        RECT 30.715 89.205 30.885 91.515 ;
        RECT 31.565 91.095 32.065 91.265 ;
        RECT 33.065 91.095 33.565 91.265 ;
        RECT 34.565 91.095 35.065 91.265 ;
        RECT 36.065 91.095 36.565 91.265 ;
        RECT 37.565 91.095 38.065 91.265 ;
        RECT 39.065 91.095 39.565 91.265 ;
        RECT 40.565 91.095 41.065 91.265 ;
        RECT 42.065 91.095 42.565 91.265 ;
        RECT 43.565 91.095 44.065 91.265 ;
        RECT 45.065 91.095 45.565 91.265 ;
        RECT 46.565 91.095 47.065 91.265 ;
        RECT 48.065 91.095 48.565 91.265 ;
        RECT 49.565 91.095 50.065 91.265 ;
        RECT 51.065 91.095 51.565 91.265 ;
        RECT 52.565 91.095 53.065 91.265 ;
        RECT 54.065 91.095 54.565 91.265 ;
        RECT 55.565 91.095 56.065 91.265 ;
        RECT 57.065 91.095 57.565 91.265 ;
        RECT 58.565 91.095 59.065 91.265 ;
        RECT 60.065 91.095 60.565 91.265 ;
        RECT 61.565 91.095 62.065 91.265 ;
        RECT 63.065 91.095 63.565 91.265 ;
        RECT 64.565 91.095 65.065 91.265 ;
        RECT 66.065 91.095 66.565 91.265 ;
        RECT 67.565 91.095 68.065 91.265 ;
        RECT 69.065 91.095 69.565 91.265 ;
        RECT 70.565 91.095 71.065 91.265 ;
        RECT 72.065 91.095 72.565 91.265 ;
        RECT 73.565 91.095 74.065 91.265 ;
        RECT 75.065 91.095 75.565 91.265 ;
        RECT 76.565 91.095 77.065 91.265 ;
        RECT 78.065 91.095 78.565 91.265 ;
        RECT 79.565 91.095 80.065 91.265 ;
        RECT 81.065 91.095 81.565 91.265 ;
        RECT 82.565 91.095 83.065 91.265 ;
        RECT 84.065 91.095 84.565 91.265 ;
        RECT 85.565 91.095 86.065 91.265 ;
        RECT 87.065 91.095 87.565 91.265 ;
        RECT 88.565 91.095 89.065 91.265 ;
        RECT 90.065 91.095 90.565 91.265 ;
        RECT 91.565 91.095 92.065 91.265 ;
        RECT 93.065 91.095 93.565 91.265 ;
        RECT 94.565 91.095 95.065 91.265 ;
        RECT 96.065 91.095 96.565 91.265 ;
        RECT 97.565 91.095 98.065 91.265 ;
        RECT 99.065 91.095 99.565 91.265 ;
        RECT 100.565 91.095 101.065 91.265 ;
        RECT 102.065 91.095 102.565 91.265 ;
        RECT 103.565 91.095 104.065 91.265 ;
        RECT 105.065 91.095 105.565 91.265 ;
        RECT 106.565 91.095 107.065 91.265 ;
        RECT 31.275 89.840 31.445 90.880 ;
        RECT 32.185 89.840 32.355 90.880 ;
        RECT 32.775 89.840 32.945 90.880 ;
        RECT 33.685 89.840 33.855 90.880 ;
        RECT 34.275 89.840 34.445 90.880 ;
        RECT 35.185 89.840 35.355 90.880 ;
        RECT 35.775 89.840 35.945 90.880 ;
        RECT 36.685 89.840 36.855 90.880 ;
        RECT 37.275 89.840 37.445 90.880 ;
        RECT 38.185 89.840 38.355 90.880 ;
        RECT 38.775 89.840 38.945 90.880 ;
        RECT 39.685 89.840 39.855 90.880 ;
        RECT 40.275 89.840 40.445 90.880 ;
        RECT 41.185 89.840 41.355 90.880 ;
        RECT 41.775 89.840 41.945 90.880 ;
        RECT 42.685 89.840 42.855 90.880 ;
        RECT 43.275 89.840 43.445 90.880 ;
        RECT 44.185 89.840 44.355 90.880 ;
        RECT 44.775 89.840 44.945 90.880 ;
        RECT 45.685 89.840 45.855 90.880 ;
        RECT 46.275 89.840 46.445 90.880 ;
        RECT 47.185 89.840 47.355 90.880 ;
        RECT 47.775 89.840 47.945 90.880 ;
        RECT 48.685 89.840 48.855 90.880 ;
        RECT 49.275 89.840 49.445 90.880 ;
        RECT 50.185 89.840 50.355 90.880 ;
        RECT 50.775 89.840 50.945 90.880 ;
        RECT 51.685 89.840 51.855 90.880 ;
        RECT 52.275 89.840 52.445 90.880 ;
        RECT 53.185 89.840 53.355 90.880 ;
        RECT 53.775 89.840 53.945 90.880 ;
        RECT 54.685 89.840 54.855 90.880 ;
        RECT 55.275 89.840 55.445 90.880 ;
        RECT 56.185 89.840 56.355 90.880 ;
        RECT 56.775 89.840 56.945 90.880 ;
        RECT 57.685 89.840 57.855 90.880 ;
        RECT 58.275 89.840 58.445 90.880 ;
        RECT 59.185 89.840 59.355 90.880 ;
        RECT 59.775 89.840 59.945 90.880 ;
        RECT 60.685 89.840 60.855 90.880 ;
        RECT 61.275 89.840 61.445 90.880 ;
        RECT 62.185 89.840 62.355 90.880 ;
        RECT 62.775 89.840 62.945 90.880 ;
        RECT 63.685 89.840 63.855 90.880 ;
        RECT 64.275 89.840 64.445 90.880 ;
        RECT 65.185 89.840 65.355 90.880 ;
        RECT 65.775 89.840 65.945 90.880 ;
        RECT 66.685 89.840 66.855 90.880 ;
        RECT 67.275 89.840 67.445 90.880 ;
        RECT 68.185 89.840 68.355 90.880 ;
        RECT 68.775 89.840 68.945 90.880 ;
        RECT 69.685 89.840 69.855 90.880 ;
        RECT 70.275 89.840 70.445 90.880 ;
        RECT 71.185 89.840 71.355 90.880 ;
        RECT 71.775 89.840 71.945 90.880 ;
        RECT 72.685 89.840 72.855 90.880 ;
        RECT 73.275 89.840 73.445 90.880 ;
        RECT 74.185 89.840 74.355 90.880 ;
        RECT 74.775 89.840 74.945 90.880 ;
        RECT 75.685 89.840 75.855 90.880 ;
        RECT 76.275 89.840 76.445 90.880 ;
        RECT 77.185 89.840 77.355 90.880 ;
        RECT 77.775 89.840 77.945 90.880 ;
        RECT 78.685 89.840 78.855 90.880 ;
        RECT 79.275 89.840 79.445 90.880 ;
        RECT 80.185 89.840 80.355 90.880 ;
        RECT 80.775 89.840 80.945 90.880 ;
        RECT 81.685 89.840 81.855 90.880 ;
        RECT 82.275 89.840 82.445 90.880 ;
        RECT 83.185 89.840 83.355 90.880 ;
        RECT 83.775 89.840 83.945 90.880 ;
        RECT 84.685 89.840 84.855 90.880 ;
        RECT 85.275 89.840 85.445 90.880 ;
        RECT 86.185 89.840 86.355 90.880 ;
        RECT 86.775 89.840 86.945 90.880 ;
        RECT 87.685 89.840 87.855 90.880 ;
        RECT 88.275 89.840 88.445 90.880 ;
        RECT 89.185 89.840 89.355 90.880 ;
        RECT 89.775 89.840 89.945 90.880 ;
        RECT 90.685 89.840 90.855 90.880 ;
        RECT 91.275 89.840 91.445 90.880 ;
        RECT 92.185 89.840 92.355 90.880 ;
        RECT 92.775 89.840 92.945 90.880 ;
        RECT 93.685 89.840 93.855 90.880 ;
        RECT 94.275 89.840 94.445 90.880 ;
        RECT 95.185 89.840 95.355 90.880 ;
        RECT 95.775 89.840 95.945 90.880 ;
        RECT 96.685 89.840 96.855 90.880 ;
        RECT 97.275 89.840 97.445 90.880 ;
        RECT 98.185 89.840 98.355 90.880 ;
        RECT 98.775 89.840 98.945 90.880 ;
        RECT 99.685 89.840 99.855 90.880 ;
        RECT 100.275 89.840 100.445 90.880 ;
        RECT 101.185 89.840 101.355 90.880 ;
        RECT 101.775 89.840 101.945 90.880 ;
        RECT 102.685 89.840 102.855 90.880 ;
        RECT 103.275 89.840 103.445 90.880 ;
        RECT 104.185 89.840 104.355 90.880 ;
        RECT 104.775 89.840 104.945 90.880 ;
        RECT 105.685 89.840 105.855 90.880 ;
        RECT 106.275 89.840 106.445 90.880 ;
        RECT 107.185 89.840 107.355 90.880 ;
        RECT 31.565 89.455 32.065 89.625 ;
        RECT 33.065 89.455 33.565 89.625 ;
        RECT 34.565 89.455 35.065 89.625 ;
        RECT 36.065 89.455 36.565 89.625 ;
        RECT 37.565 89.455 38.065 89.625 ;
        RECT 39.065 89.455 39.565 89.625 ;
        RECT 40.565 89.455 41.065 89.625 ;
        RECT 42.065 89.455 42.565 89.625 ;
        RECT 43.565 89.455 44.065 89.625 ;
        RECT 45.065 89.455 45.565 89.625 ;
        RECT 46.565 89.455 47.065 89.625 ;
        RECT 48.065 89.455 48.565 89.625 ;
        RECT 49.565 89.455 50.065 89.625 ;
        RECT 51.065 89.455 51.565 89.625 ;
        RECT 52.565 89.455 53.065 89.625 ;
        RECT 54.065 89.455 54.565 89.625 ;
        RECT 55.565 89.455 56.065 89.625 ;
        RECT 57.065 89.455 57.565 89.625 ;
        RECT 58.565 89.455 59.065 89.625 ;
        RECT 60.065 89.455 60.565 89.625 ;
        RECT 61.565 89.455 62.065 89.625 ;
        RECT 63.065 89.455 63.565 89.625 ;
        RECT 64.565 89.455 65.065 89.625 ;
        RECT 66.065 89.455 66.565 89.625 ;
        RECT 67.565 89.455 68.065 89.625 ;
        RECT 69.065 89.455 69.565 89.625 ;
        RECT 70.565 89.455 71.065 89.625 ;
        RECT 72.065 89.455 72.565 89.625 ;
        RECT 73.565 89.455 74.065 89.625 ;
        RECT 75.065 89.455 75.565 89.625 ;
        RECT 76.565 89.455 77.065 89.625 ;
        RECT 78.065 89.455 78.565 89.625 ;
        RECT 79.565 89.455 80.065 89.625 ;
        RECT 81.065 89.455 81.565 89.625 ;
        RECT 82.565 89.455 83.065 89.625 ;
        RECT 84.065 89.455 84.565 89.625 ;
        RECT 85.565 89.455 86.065 89.625 ;
        RECT 87.065 89.455 87.565 89.625 ;
        RECT 88.565 89.455 89.065 89.625 ;
        RECT 90.065 89.455 90.565 89.625 ;
        RECT 91.565 89.455 92.065 89.625 ;
        RECT 93.065 89.455 93.565 89.625 ;
        RECT 94.565 89.455 95.065 89.625 ;
        RECT 96.065 89.455 96.565 89.625 ;
        RECT 97.565 89.455 98.065 89.625 ;
        RECT 99.065 89.455 99.565 89.625 ;
        RECT 100.565 89.455 101.065 89.625 ;
        RECT 102.065 89.455 102.565 89.625 ;
        RECT 103.565 89.455 104.065 89.625 ;
        RECT 105.065 89.455 105.565 89.625 ;
        RECT 106.565 89.455 107.065 89.625 ;
        RECT 107.745 89.205 107.915 91.515 ;
        RECT 30.715 89.035 107.915 89.205 ;
        RECT 30.615 87.985 108.065 88.155 ;
        RECT 30.615 86.025 30.785 87.985 ;
        RECT 31.565 87.520 32.065 87.690 ;
        RECT 33.065 87.520 33.565 87.690 ;
        RECT 34.565 87.520 35.065 87.690 ;
        RECT 36.065 87.520 36.565 87.690 ;
        RECT 37.565 87.520 38.065 87.690 ;
        RECT 39.065 87.520 39.565 87.690 ;
        RECT 40.565 87.520 41.065 87.690 ;
        RECT 42.065 87.520 42.565 87.690 ;
        RECT 43.565 87.520 44.065 87.690 ;
        RECT 45.065 87.520 45.565 87.690 ;
        RECT 46.565 87.520 47.065 87.690 ;
        RECT 48.065 87.520 48.565 87.690 ;
        RECT 49.565 87.520 50.065 87.690 ;
        RECT 51.065 87.520 51.565 87.690 ;
        RECT 52.565 87.520 53.065 87.690 ;
        RECT 54.065 87.520 54.565 87.690 ;
        RECT 55.565 87.520 56.065 87.690 ;
        RECT 57.065 87.520 57.565 87.690 ;
        RECT 58.565 87.520 59.065 87.690 ;
        RECT 60.065 87.520 60.565 87.690 ;
        RECT 61.565 87.520 62.065 87.690 ;
        RECT 63.065 87.520 63.565 87.690 ;
        RECT 64.565 87.520 65.065 87.690 ;
        RECT 66.065 87.520 66.565 87.690 ;
        RECT 67.565 87.520 68.065 87.690 ;
        RECT 69.065 87.520 69.565 87.690 ;
        RECT 70.565 87.520 71.065 87.690 ;
        RECT 72.065 87.520 72.565 87.690 ;
        RECT 73.565 87.520 74.065 87.690 ;
        RECT 75.065 87.520 75.565 87.690 ;
        RECT 76.565 87.520 77.065 87.690 ;
        RECT 78.065 87.520 78.565 87.690 ;
        RECT 79.565 87.520 80.065 87.690 ;
        RECT 81.065 87.520 81.565 87.690 ;
        RECT 82.565 87.520 83.065 87.690 ;
        RECT 84.065 87.520 84.565 87.690 ;
        RECT 85.565 87.520 86.065 87.690 ;
        RECT 87.065 87.520 87.565 87.690 ;
        RECT 88.565 87.520 89.065 87.690 ;
        RECT 90.065 87.520 90.565 87.690 ;
        RECT 91.565 87.520 92.065 87.690 ;
        RECT 93.065 87.520 93.565 87.690 ;
        RECT 94.565 87.520 95.065 87.690 ;
        RECT 96.065 87.520 96.565 87.690 ;
        RECT 97.565 87.520 98.065 87.690 ;
        RECT 99.065 87.520 99.565 87.690 ;
        RECT 100.565 87.520 101.065 87.690 ;
        RECT 102.065 87.520 102.565 87.690 ;
        RECT 103.565 87.520 104.065 87.690 ;
        RECT 105.065 87.520 105.565 87.690 ;
        RECT 106.565 87.520 107.065 87.690 ;
        RECT 31.275 86.660 31.445 87.350 ;
        RECT 32.185 86.660 32.355 87.350 ;
        RECT 32.775 86.660 32.945 87.350 ;
        RECT 33.685 86.660 33.855 87.350 ;
        RECT 34.275 86.660 34.445 87.350 ;
        RECT 35.185 86.660 35.355 87.350 ;
        RECT 35.775 86.660 35.945 87.350 ;
        RECT 36.685 86.660 36.855 87.350 ;
        RECT 37.275 86.660 37.445 87.350 ;
        RECT 38.185 86.660 38.355 87.350 ;
        RECT 38.775 86.660 38.945 87.350 ;
        RECT 39.685 86.660 39.855 87.350 ;
        RECT 40.275 86.660 40.445 87.350 ;
        RECT 41.185 86.660 41.355 87.350 ;
        RECT 41.775 86.660 41.945 87.350 ;
        RECT 42.685 86.660 42.855 87.350 ;
        RECT 43.275 86.660 43.445 87.350 ;
        RECT 44.185 86.660 44.355 87.350 ;
        RECT 44.775 86.660 44.945 87.350 ;
        RECT 45.685 86.660 45.855 87.350 ;
        RECT 46.275 86.660 46.445 87.350 ;
        RECT 47.185 86.660 47.355 87.350 ;
        RECT 47.775 86.660 47.945 87.350 ;
        RECT 48.685 86.660 48.855 87.350 ;
        RECT 49.275 86.660 49.445 87.350 ;
        RECT 50.185 86.660 50.355 87.350 ;
        RECT 50.775 86.660 50.945 87.350 ;
        RECT 51.685 86.660 51.855 87.350 ;
        RECT 52.275 86.660 52.445 87.350 ;
        RECT 53.185 86.660 53.355 87.350 ;
        RECT 53.775 86.660 53.945 87.350 ;
        RECT 54.685 86.660 54.855 87.350 ;
        RECT 55.275 86.660 55.445 87.350 ;
        RECT 56.185 86.660 56.355 87.350 ;
        RECT 56.775 86.660 56.945 87.350 ;
        RECT 57.685 86.660 57.855 87.350 ;
        RECT 58.275 86.660 58.445 87.350 ;
        RECT 59.185 86.660 59.355 87.350 ;
        RECT 59.775 86.660 59.945 87.350 ;
        RECT 60.685 86.660 60.855 87.350 ;
        RECT 61.275 86.660 61.445 87.350 ;
        RECT 62.185 86.660 62.355 87.350 ;
        RECT 62.775 86.660 62.945 87.350 ;
        RECT 63.685 86.660 63.855 87.350 ;
        RECT 64.275 86.660 64.445 87.350 ;
        RECT 65.185 86.660 65.355 87.350 ;
        RECT 65.775 86.660 65.945 87.350 ;
        RECT 66.685 86.660 66.855 87.350 ;
        RECT 67.275 86.660 67.445 87.350 ;
        RECT 68.185 86.660 68.355 87.350 ;
        RECT 68.775 86.660 68.945 87.350 ;
        RECT 69.685 86.660 69.855 87.350 ;
        RECT 70.275 86.660 70.445 87.350 ;
        RECT 71.185 86.660 71.355 87.350 ;
        RECT 71.775 86.660 71.945 87.350 ;
        RECT 72.685 86.660 72.855 87.350 ;
        RECT 73.275 86.660 73.445 87.350 ;
        RECT 74.185 86.660 74.355 87.350 ;
        RECT 74.775 86.660 74.945 87.350 ;
        RECT 75.685 86.660 75.855 87.350 ;
        RECT 76.275 86.660 76.445 87.350 ;
        RECT 77.185 86.660 77.355 87.350 ;
        RECT 77.775 86.660 77.945 87.350 ;
        RECT 78.685 86.660 78.855 87.350 ;
        RECT 79.275 86.660 79.445 87.350 ;
        RECT 80.185 86.660 80.355 87.350 ;
        RECT 80.775 86.660 80.945 87.350 ;
        RECT 81.685 86.660 81.855 87.350 ;
        RECT 82.275 86.660 82.445 87.350 ;
        RECT 83.185 86.660 83.355 87.350 ;
        RECT 83.775 86.660 83.945 87.350 ;
        RECT 84.685 86.660 84.855 87.350 ;
        RECT 85.275 86.660 85.445 87.350 ;
        RECT 86.185 86.660 86.355 87.350 ;
        RECT 86.775 86.660 86.945 87.350 ;
        RECT 87.685 86.660 87.855 87.350 ;
        RECT 88.275 86.660 88.445 87.350 ;
        RECT 89.185 86.660 89.355 87.350 ;
        RECT 89.775 86.660 89.945 87.350 ;
        RECT 90.685 86.660 90.855 87.350 ;
        RECT 91.275 86.660 91.445 87.350 ;
        RECT 92.185 86.660 92.355 87.350 ;
        RECT 92.775 86.660 92.945 87.350 ;
        RECT 93.685 86.660 93.855 87.350 ;
        RECT 94.275 86.660 94.445 87.350 ;
        RECT 95.185 86.660 95.355 87.350 ;
        RECT 95.775 86.660 95.945 87.350 ;
        RECT 96.685 86.660 96.855 87.350 ;
        RECT 97.275 86.660 97.445 87.350 ;
        RECT 98.185 86.660 98.355 87.350 ;
        RECT 98.775 86.660 98.945 87.350 ;
        RECT 99.685 86.660 99.855 87.350 ;
        RECT 100.275 86.660 100.445 87.350 ;
        RECT 101.185 86.660 101.355 87.350 ;
        RECT 101.775 86.660 101.945 87.350 ;
        RECT 102.685 86.660 102.855 87.350 ;
        RECT 103.275 86.660 103.445 87.350 ;
        RECT 104.185 86.660 104.355 87.350 ;
        RECT 104.775 86.660 104.945 87.350 ;
        RECT 105.685 86.660 105.855 87.350 ;
        RECT 106.275 86.660 106.445 87.350 ;
        RECT 107.185 86.660 107.355 87.350 ;
        RECT 31.565 86.320 32.065 86.490 ;
        RECT 33.065 86.320 33.565 86.490 ;
        RECT 34.565 86.320 35.065 86.490 ;
        RECT 36.065 86.320 36.565 86.490 ;
        RECT 37.565 86.320 38.065 86.490 ;
        RECT 39.065 86.320 39.565 86.490 ;
        RECT 40.565 86.320 41.065 86.490 ;
        RECT 42.065 86.320 42.565 86.490 ;
        RECT 43.565 86.320 44.065 86.490 ;
        RECT 45.065 86.320 45.565 86.490 ;
        RECT 46.565 86.320 47.065 86.490 ;
        RECT 48.065 86.320 48.565 86.490 ;
        RECT 49.565 86.320 50.065 86.490 ;
        RECT 51.065 86.320 51.565 86.490 ;
        RECT 52.565 86.320 53.065 86.490 ;
        RECT 54.065 86.320 54.565 86.490 ;
        RECT 55.565 86.320 56.065 86.490 ;
        RECT 57.065 86.320 57.565 86.490 ;
        RECT 58.565 86.320 59.065 86.490 ;
        RECT 60.065 86.320 60.565 86.490 ;
        RECT 61.565 86.320 62.065 86.490 ;
        RECT 63.065 86.320 63.565 86.490 ;
        RECT 64.565 86.320 65.065 86.490 ;
        RECT 66.065 86.320 66.565 86.490 ;
        RECT 67.565 86.320 68.065 86.490 ;
        RECT 69.065 86.320 69.565 86.490 ;
        RECT 70.565 86.320 71.065 86.490 ;
        RECT 72.065 86.320 72.565 86.490 ;
        RECT 73.565 86.320 74.065 86.490 ;
        RECT 75.065 86.320 75.565 86.490 ;
        RECT 76.565 86.320 77.065 86.490 ;
        RECT 78.065 86.320 78.565 86.490 ;
        RECT 79.565 86.320 80.065 86.490 ;
        RECT 81.065 86.320 81.565 86.490 ;
        RECT 82.565 86.320 83.065 86.490 ;
        RECT 84.065 86.320 84.565 86.490 ;
        RECT 85.565 86.320 86.065 86.490 ;
        RECT 87.065 86.320 87.565 86.490 ;
        RECT 88.565 86.320 89.065 86.490 ;
        RECT 90.065 86.320 90.565 86.490 ;
        RECT 91.565 86.320 92.065 86.490 ;
        RECT 93.065 86.320 93.565 86.490 ;
        RECT 94.565 86.320 95.065 86.490 ;
        RECT 96.065 86.320 96.565 86.490 ;
        RECT 97.565 86.320 98.065 86.490 ;
        RECT 99.065 86.320 99.565 86.490 ;
        RECT 100.565 86.320 101.065 86.490 ;
        RECT 102.065 86.320 102.565 86.490 ;
        RECT 103.565 86.320 104.065 86.490 ;
        RECT 105.065 86.320 105.565 86.490 ;
        RECT 106.565 86.320 107.065 86.490 ;
        RECT 107.895 86.025 108.065 87.985 ;
        RECT 30.615 85.855 108.065 86.025 ;
        RECT 36.380 78.680 39.030 78.850 ;
        RECT 36.380 64.820 36.550 78.680 ;
        RECT 37.185 78.120 38.225 78.290 ;
        RECT 36.800 77.500 36.970 78.000 ;
        RECT 38.440 77.500 38.610 78.000 ;
        RECT 37.185 77.210 38.225 77.380 ;
        RECT 37.185 76.620 38.225 76.790 ;
        RECT 36.800 76.000 36.970 76.500 ;
        RECT 38.440 76.000 38.610 76.500 ;
        RECT 37.185 75.710 38.225 75.880 ;
        RECT 37.185 75.120 38.225 75.290 ;
        RECT 36.800 74.500 36.970 75.000 ;
        RECT 38.440 74.500 38.610 75.000 ;
        RECT 37.185 74.210 38.225 74.380 ;
        RECT 37.185 73.620 38.225 73.790 ;
        RECT 36.800 73.000 36.970 73.500 ;
        RECT 38.440 73.000 38.610 73.500 ;
        RECT 37.185 72.710 38.225 72.880 ;
        RECT 37.185 72.120 38.225 72.290 ;
        RECT 36.800 71.500 36.970 72.000 ;
        RECT 38.440 71.500 38.610 72.000 ;
        RECT 37.185 71.210 38.225 71.380 ;
        RECT 37.185 70.620 38.225 70.790 ;
        RECT 36.800 70.000 36.970 70.500 ;
        RECT 38.440 70.000 38.610 70.500 ;
        RECT 37.185 69.710 38.225 69.880 ;
        RECT 37.185 69.120 38.225 69.290 ;
        RECT 36.800 68.500 36.970 69.000 ;
        RECT 38.440 68.500 38.610 69.000 ;
        RECT 37.185 68.210 38.225 68.380 ;
        RECT 37.185 67.620 38.225 67.790 ;
        RECT 36.800 67.000 36.970 67.500 ;
        RECT 38.440 67.000 38.610 67.500 ;
        RECT 37.185 66.710 38.225 66.880 ;
        RECT 37.185 66.120 38.225 66.290 ;
        RECT 36.800 65.500 36.970 66.000 ;
        RECT 38.440 65.500 38.610 66.000 ;
        RECT 37.185 65.210 38.225 65.380 ;
        RECT 38.860 64.820 39.030 78.680 ;
        RECT 36.380 64.650 39.030 64.820 ;
        RECT 39.910 78.830 42.210 79.000 ;
        RECT 39.910 64.720 40.080 78.830 ;
        RECT 40.715 78.120 41.405 78.290 ;
        RECT 40.375 77.500 40.545 78.000 ;
        RECT 41.575 77.500 41.745 78.000 ;
        RECT 40.715 77.210 41.405 77.380 ;
        RECT 40.715 76.620 41.405 76.790 ;
        RECT 40.375 76.000 40.545 76.500 ;
        RECT 41.575 76.000 41.745 76.500 ;
        RECT 40.715 75.710 41.405 75.880 ;
        RECT 40.715 75.120 41.405 75.290 ;
        RECT 40.375 74.500 40.545 75.000 ;
        RECT 41.575 74.500 41.745 75.000 ;
        RECT 40.715 74.210 41.405 74.380 ;
        RECT 40.715 73.620 41.405 73.790 ;
        RECT 40.375 73.000 40.545 73.500 ;
        RECT 41.575 73.000 41.745 73.500 ;
        RECT 40.715 72.710 41.405 72.880 ;
        RECT 40.715 72.120 41.405 72.290 ;
        RECT 40.375 71.500 40.545 72.000 ;
        RECT 41.575 71.500 41.745 72.000 ;
        RECT 40.715 71.210 41.405 71.380 ;
        RECT 40.715 70.620 41.405 70.790 ;
        RECT 40.375 70.000 40.545 70.500 ;
        RECT 41.575 70.000 41.745 70.500 ;
        RECT 40.715 69.710 41.405 69.880 ;
        RECT 40.715 69.120 41.405 69.290 ;
        RECT 40.375 68.500 40.545 69.000 ;
        RECT 41.575 68.500 41.745 69.000 ;
        RECT 40.715 68.210 41.405 68.380 ;
        RECT 40.715 67.620 41.405 67.790 ;
        RECT 40.375 67.000 40.545 67.500 ;
        RECT 41.575 67.000 41.745 67.500 ;
        RECT 40.715 66.710 41.405 66.880 ;
        RECT 40.715 66.120 41.405 66.290 ;
        RECT 40.375 65.500 40.545 66.000 ;
        RECT 41.575 65.500 41.745 66.000 ;
        RECT 40.715 65.210 41.405 65.380 ;
        RECT 42.040 64.720 42.210 78.830 ;
        RECT 39.910 64.550 42.210 64.720 ;
        RECT 43.090 78.680 45.740 78.850 ;
        RECT 43.090 64.820 43.260 78.680 ;
        RECT 43.895 78.120 44.935 78.290 ;
        RECT 43.510 77.500 43.680 78.000 ;
        RECT 45.150 77.500 45.320 78.000 ;
        RECT 43.895 77.210 44.935 77.380 ;
        RECT 43.895 76.620 44.935 76.790 ;
        RECT 43.510 76.000 43.680 76.500 ;
        RECT 45.150 76.000 45.320 76.500 ;
        RECT 43.895 75.710 44.935 75.880 ;
        RECT 43.895 75.120 44.935 75.290 ;
        RECT 43.510 74.500 43.680 75.000 ;
        RECT 45.150 74.500 45.320 75.000 ;
        RECT 43.895 74.210 44.935 74.380 ;
        RECT 43.895 73.620 44.935 73.790 ;
        RECT 43.510 73.000 43.680 73.500 ;
        RECT 45.150 73.000 45.320 73.500 ;
        RECT 43.895 72.710 44.935 72.880 ;
        RECT 43.895 72.120 44.935 72.290 ;
        RECT 43.510 71.500 43.680 72.000 ;
        RECT 45.150 71.500 45.320 72.000 ;
        RECT 43.895 71.210 44.935 71.380 ;
        RECT 43.895 70.620 44.935 70.790 ;
        RECT 43.510 70.000 43.680 70.500 ;
        RECT 45.150 70.000 45.320 70.500 ;
        RECT 43.895 69.710 44.935 69.880 ;
        RECT 43.895 69.120 44.935 69.290 ;
        RECT 43.510 68.500 43.680 69.000 ;
        RECT 45.150 68.500 45.320 69.000 ;
        RECT 43.895 68.210 44.935 68.380 ;
        RECT 43.895 67.620 44.935 67.790 ;
        RECT 43.510 67.000 43.680 67.500 ;
        RECT 45.150 67.000 45.320 67.500 ;
        RECT 43.895 66.710 44.935 66.880 ;
        RECT 43.895 66.120 44.935 66.290 ;
        RECT 43.510 65.500 43.680 66.000 ;
        RECT 45.150 65.500 45.320 66.000 ;
        RECT 43.895 65.210 44.935 65.380 ;
        RECT 45.570 64.820 45.740 78.680 ;
        RECT 43.090 64.650 45.740 64.820 ;
        RECT 46.620 78.830 48.920 79.000 ;
        RECT 46.620 64.720 46.790 78.830 ;
        RECT 47.425 78.120 48.115 78.290 ;
        RECT 47.085 77.500 47.255 78.000 ;
        RECT 48.285 77.500 48.455 78.000 ;
        RECT 47.425 77.210 48.115 77.380 ;
        RECT 47.425 76.620 48.115 76.790 ;
        RECT 47.085 76.000 47.255 76.500 ;
        RECT 48.285 76.000 48.455 76.500 ;
        RECT 47.425 75.710 48.115 75.880 ;
        RECT 47.425 75.120 48.115 75.290 ;
        RECT 47.085 74.500 47.255 75.000 ;
        RECT 48.285 74.500 48.455 75.000 ;
        RECT 47.425 74.210 48.115 74.380 ;
        RECT 47.425 73.620 48.115 73.790 ;
        RECT 47.085 73.000 47.255 73.500 ;
        RECT 48.285 73.000 48.455 73.500 ;
        RECT 47.425 72.710 48.115 72.880 ;
        RECT 47.425 72.120 48.115 72.290 ;
        RECT 47.085 71.500 47.255 72.000 ;
        RECT 48.285 71.500 48.455 72.000 ;
        RECT 47.425 71.210 48.115 71.380 ;
        RECT 47.425 70.620 48.115 70.790 ;
        RECT 47.085 70.000 47.255 70.500 ;
        RECT 48.285 70.000 48.455 70.500 ;
        RECT 47.425 69.710 48.115 69.880 ;
        RECT 47.425 69.120 48.115 69.290 ;
        RECT 47.085 68.500 47.255 69.000 ;
        RECT 48.285 68.500 48.455 69.000 ;
        RECT 47.425 68.210 48.115 68.380 ;
        RECT 47.425 67.620 48.115 67.790 ;
        RECT 47.085 67.000 47.255 67.500 ;
        RECT 48.285 67.000 48.455 67.500 ;
        RECT 47.425 66.710 48.115 66.880 ;
        RECT 47.425 66.120 48.115 66.290 ;
        RECT 47.085 65.500 47.255 66.000 ;
        RECT 48.285 65.500 48.455 66.000 ;
        RECT 47.425 65.210 48.115 65.380 ;
        RECT 48.750 64.720 48.920 78.830 ;
        RECT 46.620 64.550 48.920 64.720 ;
        RECT 49.800 78.680 52.450 78.850 ;
        RECT 49.800 64.820 49.970 78.680 ;
        RECT 50.605 78.120 51.645 78.290 ;
        RECT 50.220 77.500 50.390 78.000 ;
        RECT 51.860 77.500 52.030 78.000 ;
        RECT 50.605 77.210 51.645 77.380 ;
        RECT 50.605 76.620 51.645 76.790 ;
        RECT 50.220 76.000 50.390 76.500 ;
        RECT 51.860 76.000 52.030 76.500 ;
        RECT 50.605 75.710 51.645 75.880 ;
        RECT 50.605 75.120 51.645 75.290 ;
        RECT 50.220 74.500 50.390 75.000 ;
        RECT 51.860 74.500 52.030 75.000 ;
        RECT 50.605 74.210 51.645 74.380 ;
        RECT 50.605 73.620 51.645 73.790 ;
        RECT 50.220 73.000 50.390 73.500 ;
        RECT 51.860 73.000 52.030 73.500 ;
        RECT 50.605 72.710 51.645 72.880 ;
        RECT 50.605 72.120 51.645 72.290 ;
        RECT 50.220 71.500 50.390 72.000 ;
        RECT 51.860 71.500 52.030 72.000 ;
        RECT 50.605 71.210 51.645 71.380 ;
        RECT 50.605 70.620 51.645 70.790 ;
        RECT 50.220 70.000 50.390 70.500 ;
        RECT 51.860 70.000 52.030 70.500 ;
        RECT 50.605 69.710 51.645 69.880 ;
        RECT 50.605 69.120 51.645 69.290 ;
        RECT 50.220 68.500 50.390 69.000 ;
        RECT 51.860 68.500 52.030 69.000 ;
        RECT 50.605 68.210 51.645 68.380 ;
        RECT 50.605 67.620 51.645 67.790 ;
        RECT 50.220 67.000 50.390 67.500 ;
        RECT 51.860 67.000 52.030 67.500 ;
        RECT 50.605 66.710 51.645 66.880 ;
        RECT 50.605 66.120 51.645 66.290 ;
        RECT 50.220 65.500 50.390 66.000 ;
        RECT 51.860 65.500 52.030 66.000 ;
        RECT 50.605 65.210 51.645 65.380 ;
        RECT 52.280 64.820 52.450 78.680 ;
        RECT 49.800 64.650 52.450 64.820 ;
        RECT 53.330 78.830 55.630 79.000 ;
        RECT 53.330 64.720 53.500 78.830 ;
        RECT 54.135 78.120 54.825 78.290 ;
        RECT 53.795 77.500 53.965 78.000 ;
        RECT 54.995 77.500 55.165 78.000 ;
        RECT 54.135 77.210 54.825 77.380 ;
        RECT 54.135 76.620 54.825 76.790 ;
        RECT 53.795 76.000 53.965 76.500 ;
        RECT 54.995 76.000 55.165 76.500 ;
        RECT 54.135 75.710 54.825 75.880 ;
        RECT 54.135 75.120 54.825 75.290 ;
        RECT 53.795 74.500 53.965 75.000 ;
        RECT 54.995 74.500 55.165 75.000 ;
        RECT 54.135 74.210 54.825 74.380 ;
        RECT 54.135 73.620 54.825 73.790 ;
        RECT 53.795 73.000 53.965 73.500 ;
        RECT 54.995 73.000 55.165 73.500 ;
        RECT 54.135 72.710 54.825 72.880 ;
        RECT 54.135 72.120 54.825 72.290 ;
        RECT 53.795 71.500 53.965 72.000 ;
        RECT 54.995 71.500 55.165 72.000 ;
        RECT 54.135 71.210 54.825 71.380 ;
        RECT 54.135 70.620 54.825 70.790 ;
        RECT 53.795 70.000 53.965 70.500 ;
        RECT 54.995 70.000 55.165 70.500 ;
        RECT 54.135 69.710 54.825 69.880 ;
        RECT 54.135 69.120 54.825 69.290 ;
        RECT 53.795 68.500 53.965 69.000 ;
        RECT 54.995 68.500 55.165 69.000 ;
        RECT 54.135 68.210 54.825 68.380 ;
        RECT 54.135 67.620 54.825 67.790 ;
        RECT 53.795 67.000 53.965 67.500 ;
        RECT 54.995 67.000 55.165 67.500 ;
        RECT 54.135 66.710 54.825 66.880 ;
        RECT 54.135 66.120 54.825 66.290 ;
        RECT 53.795 65.500 53.965 66.000 ;
        RECT 54.995 65.500 55.165 66.000 ;
        RECT 54.135 65.210 54.825 65.380 ;
        RECT 55.460 64.720 55.630 78.830 ;
        RECT 53.330 64.550 55.630 64.720 ;
        RECT 56.510 78.680 59.160 78.850 ;
        RECT 56.510 64.820 56.680 78.680 ;
        RECT 57.315 78.120 58.355 78.290 ;
        RECT 56.930 77.500 57.100 78.000 ;
        RECT 58.570 77.500 58.740 78.000 ;
        RECT 57.315 77.210 58.355 77.380 ;
        RECT 57.315 76.620 58.355 76.790 ;
        RECT 56.930 76.000 57.100 76.500 ;
        RECT 58.570 76.000 58.740 76.500 ;
        RECT 57.315 75.710 58.355 75.880 ;
        RECT 57.315 75.120 58.355 75.290 ;
        RECT 56.930 74.500 57.100 75.000 ;
        RECT 58.570 74.500 58.740 75.000 ;
        RECT 57.315 74.210 58.355 74.380 ;
        RECT 57.315 73.620 58.355 73.790 ;
        RECT 56.930 73.000 57.100 73.500 ;
        RECT 58.570 73.000 58.740 73.500 ;
        RECT 57.315 72.710 58.355 72.880 ;
        RECT 57.315 72.120 58.355 72.290 ;
        RECT 56.930 71.500 57.100 72.000 ;
        RECT 58.570 71.500 58.740 72.000 ;
        RECT 57.315 71.210 58.355 71.380 ;
        RECT 57.315 70.620 58.355 70.790 ;
        RECT 56.930 70.000 57.100 70.500 ;
        RECT 58.570 70.000 58.740 70.500 ;
        RECT 57.315 69.710 58.355 69.880 ;
        RECT 57.315 69.120 58.355 69.290 ;
        RECT 56.930 68.500 57.100 69.000 ;
        RECT 58.570 68.500 58.740 69.000 ;
        RECT 57.315 68.210 58.355 68.380 ;
        RECT 57.315 67.620 58.355 67.790 ;
        RECT 56.930 67.000 57.100 67.500 ;
        RECT 58.570 67.000 58.740 67.500 ;
        RECT 57.315 66.710 58.355 66.880 ;
        RECT 57.315 66.120 58.355 66.290 ;
        RECT 56.930 65.500 57.100 66.000 ;
        RECT 58.570 65.500 58.740 66.000 ;
        RECT 57.315 65.210 58.355 65.380 ;
        RECT 58.990 64.820 59.160 78.680 ;
        RECT 56.510 64.650 59.160 64.820 ;
        RECT 60.040 78.830 62.340 79.000 ;
        RECT 60.040 64.720 60.210 78.830 ;
        RECT 60.845 78.120 61.535 78.290 ;
        RECT 60.505 77.500 60.675 78.000 ;
        RECT 61.705 77.500 61.875 78.000 ;
        RECT 60.845 77.210 61.535 77.380 ;
        RECT 60.845 76.620 61.535 76.790 ;
        RECT 60.505 76.000 60.675 76.500 ;
        RECT 61.705 76.000 61.875 76.500 ;
        RECT 60.845 75.710 61.535 75.880 ;
        RECT 60.845 75.120 61.535 75.290 ;
        RECT 60.505 74.500 60.675 75.000 ;
        RECT 61.705 74.500 61.875 75.000 ;
        RECT 60.845 74.210 61.535 74.380 ;
        RECT 60.845 73.620 61.535 73.790 ;
        RECT 60.505 73.000 60.675 73.500 ;
        RECT 61.705 73.000 61.875 73.500 ;
        RECT 60.845 72.710 61.535 72.880 ;
        RECT 60.845 72.120 61.535 72.290 ;
        RECT 60.505 71.500 60.675 72.000 ;
        RECT 61.705 71.500 61.875 72.000 ;
        RECT 60.845 71.210 61.535 71.380 ;
        RECT 60.845 70.620 61.535 70.790 ;
        RECT 60.505 70.000 60.675 70.500 ;
        RECT 61.705 70.000 61.875 70.500 ;
        RECT 60.845 69.710 61.535 69.880 ;
        RECT 60.845 69.120 61.535 69.290 ;
        RECT 60.505 68.500 60.675 69.000 ;
        RECT 61.705 68.500 61.875 69.000 ;
        RECT 60.845 68.210 61.535 68.380 ;
        RECT 60.845 67.620 61.535 67.790 ;
        RECT 60.505 67.000 60.675 67.500 ;
        RECT 61.705 67.000 61.875 67.500 ;
        RECT 60.845 66.710 61.535 66.880 ;
        RECT 60.845 66.120 61.535 66.290 ;
        RECT 60.505 65.500 60.675 66.000 ;
        RECT 61.705 65.500 61.875 66.000 ;
        RECT 60.845 65.210 61.535 65.380 ;
        RECT 62.170 64.720 62.340 78.830 ;
        RECT 60.040 64.550 62.340 64.720 ;
        RECT 63.220 78.680 65.870 78.850 ;
        RECT 63.220 64.820 63.390 78.680 ;
        RECT 64.025 78.120 65.065 78.290 ;
        RECT 63.640 77.500 63.810 78.000 ;
        RECT 65.280 77.500 65.450 78.000 ;
        RECT 64.025 77.210 65.065 77.380 ;
        RECT 64.025 76.620 65.065 76.790 ;
        RECT 63.640 76.000 63.810 76.500 ;
        RECT 65.280 76.000 65.450 76.500 ;
        RECT 64.025 75.710 65.065 75.880 ;
        RECT 64.025 75.120 65.065 75.290 ;
        RECT 63.640 74.500 63.810 75.000 ;
        RECT 65.280 74.500 65.450 75.000 ;
        RECT 64.025 74.210 65.065 74.380 ;
        RECT 64.025 73.620 65.065 73.790 ;
        RECT 63.640 73.000 63.810 73.500 ;
        RECT 65.280 73.000 65.450 73.500 ;
        RECT 64.025 72.710 65.065 72.880 ;
        RECT 64.025 72.120 65.065 72.290 ;
        RECT 63.640 71.500 63.810 72.000 ;
        RECT 65.280 71.500 65.450 72.000 ;
        RECT 64.025 71.210 65.065 71.380 ;
        RECT 64.025 70.620 65.065 70.790 ;
        RECT 63.640 70.000 63.810 70.500 ;
        RECT 65.280 70.000 65.450 70.500 ;
        RECT 64.025 69.710 65.065 69.880 ;
        RECT 64.025 69.120 65.065 69.290 ;
        RECT 63.640 68.500 63.810 69.000 ;
        RECT 65.280 68.500 65.450 69.000 ;
        RECT 64.025 68.210 65.065 68.380 ;
        RECT 64.025 67.620 65.065 67.790 ;
        RECT 63.640 67.000 63.810 67.500 ;
        RECT 65.280 67.000 65.450 67.500 ;
        RECT 64.025 66.710 65.065 66.880 ;
        RECT 64.025 66.120 65.065 66.290 ;
        RECT 63.640 65.500 63.810 66.000 ;
        RECT 65.280 65.500 65.450 66.000 ;
        RECT 64.025 65.210 65.065 65.380 ;
        RECT 65.700 64.820 65.870 78.680 ;
        RECT 63.220 64.650 65.870 64.820 ;
        RECT 66.750 78.830 69.050 79.000 ;
        RECT 66.750 64.720 66.920 78.830 ;
        RECT 67.555 78.120 68.245 78.290 ;
        RECT 67.215 77.500 67.385 78.000 ;
        RECT 68.415 77.500 68.585 78.000 ;
        RECT 67.555 77.210 68.245 77.380 ;
        RECT 67.555 76.620 68.245 76.790 ;
        RECT 67.215 76.000 67.385 76.500 ;
        RECT 68.415 76.000 68.585 76.500 ;
        RECT 67.555 75.710 68.245 75.880 ;
        RECT 67.555 75.120 68.245 75.290 ;
        RECT 67.215 74.500 67.385 75.000 ;
        RECT 68.415 74.500 68.585 75.000 ;
        RECT 67.555 74.210 68.245 74.380 ;
        RECT 67.555 73.620 68.245 73.790 ;
        RECT 67.215 73.000 67.385 73.500 ;
        RECT 68.415 73.000 68.585 73.500 ;
        RECT 67.555 72.710 68.245 72.880 ;
        RECT 67.555 72.120 68.245 72.290 ;
        RECT 67.215 71.500 67.385 72.000 ;
        RECT 68.415 71.500 68.585 72.000 ;
        RECT 67.555 71.210 68.245 71.380 ;
        RECT 67.555 70.620 68.245 70.790 ;
        RECT 67.215 70.000 67.385 70.500 ;
        RECT 68.415 70.000 68.585 70.500 ;
        RECT 67.555 69.710 68.245 69.880 ;
        RECT 67.555 69.120 68.245 69.290 ;
        RECT 67.215 68.500 67.385 69.000 ;
        RECT 68.415 68.500 68.585 69.000 ;
        RECT 67.555 68.210 68.245 68.380 ;
        RECT 67.555 67.620 68.245 67.790 ;
        RECT 67.215 67.000 67.385 67.500 ;
        RECT 68.415 67.000 68.585 67.500 ;
        RECT 67.555 66.710 68.245 66.880 ;
        RECT 67.555 66.120 68.245 66.290 ;
        RECT 67.215 65.500 67.385 66.000 ;
        RECT 68.415 65.500 68.585 66.000 ;
        RECT 67.555 65.210 68.245 65.380 ;
        RECT 68.880 64.720 69.050 78.830 ;
        RECT 66.750 64.550 69.050 64.720 ;
        RECT 69.930 78.680 72.580 78.850 ;
        RECT 69.930 64.820 70.100 78.680 ;
        RECT 70.735 78.120 71.775 78.290 ;
        RECT 70.350 77.500 70.520 78.000 ;
        RECT 71.990 77.500 72.160 78.000 ;
        RECT 70.735 77.210 71.775 77.380 ;
        RECT 70.735 76.620 71.775 76.790 ;
        RECT 70.350 76.000 70.520 76.500 ;
        RECT 71.990 76.000 72.160 76.500 ;
        RECT 70.735 75.710 71.775 75.880 ;
        RECT 70.735 75.120 71.775 75.290 ;
        RECT 70.350 74.500 70.520 75.000 ;
        RECT 71.990 74.500 72.160 75.000 ;
        RECT 70.735 74.210 71.775 74.380 ;
        RECT 70.735 73.620 71.775 73.790 ;
        RECT 70.350 73.000 70.520 73.500 ;
        RECT 71.990 73.000 72.160 73.500 ;
        RECT 70.735 72.710 71.775 72.880 ;
        RECT 70.735 72.120 71.775 72.290 ;
        RECT 70.350 71.500 70.520 72.000 ;
        RECT 71.990 71.500 72.160 72.000 ;
        RECT 70.735 71.210 71.775 71.380 ;
        RECT 70.735 70.620 71.775 70.790 ;
        RECT 70.350 70.000 70.520 70.500 ;
        RECT 71.990 70.000 72.160 70.500 ;
        RECT 70.735 69.710 71.775 69.880 ;
        RECT 70.735 69.120 71.775 69.290 ;
        RECT 70.350 68.500 70.520 69.000 ;
        RECT 71.990 68.500 72.160 69.000 ;
        RECT 70.735 68.210 71.775 68.380 ;
        RECT 70.735 67.620 71.775 67.790 ;
        RECT 70.350 67.000 70.520 67.500 ;
        RECT 71.990 67.000 72.160 67.500 ;
        RECT 70.735 66.710 71.775 66.880 ;
        RECT 70.735 66.120 71.775 66.290 ;
        RECT 70.350 65.500 70.520 66.000 ;
        RECT 71.990 65.500 72.160 66.000 ;
        RECT 70.735 65.210 71.775 65.380 ;
        RECT 72.410 64.820 72.580 78.680 ;
        RECT 69.930 64.650 72.580 64.820 ;
        RECT 73.460 78.830 75.760 79.000 ;
        RECT 73.460 64.720 73.630 78.830 ;
        RECT 74.265 78.120 74.955 78.290 ;
        RECT 73.925 77.500 74.095 78.000 ;
        RECT 75.125 77.500 75.295 78.000 ;
        RECT 74.265 77.210 74.955 77.380 ;
        RECT 74.265 76.620 74.955 76.790 ;
        RECT 73.925 76.000 74.095 76.500 ;
        RECT 75.125 76.000 75.295 76.500 ;
        RECT 74.265 75.710 74.955 75.880 ;
        RECT 74.265 75.120 74.955 75.290 ;
        RECT 73.925 74.500 74.095 75.000 ;
        RECT 75.125 74.500 75.295 75.000 ;
        RECT 74.265 74.210 74.955 74.380 ;
        RECT 74.265 73.620 74.955 73.790 ;
        RECT 73.925 73.000 74.095 73.500 ;
        RECT 75.125 73.000 75.295 73.500 ;
        RECT 74.265 72.710 74.955 72.880 ;
        RECT 74.265 72.120 74.955 72.290 ;
        RECT 73.925 71.500 74.095 72.000 ;
        RECT 75.125 71.500 75.295 72.000 ;
        RECT 74.265 71.210 74.955 71.380 ;
        RECT 74.265 70.620 74.955 70.790 ;
        RECT 73.925 70.000 74.095 70.500 ;
        RECT 75.125 70.000 75.295 70.500 ;
        RECT 74.265 69.710 74.955 69.880 ;
        RECT 74.265 69.120 74.955 69.290 ;
        RECT 73.925 68.500 74.095 69.000 ;
        RECT 75.125 68.500 75.295 69.000 ;
        RECT 74.265 68.210 74.955 68.380 ;
        RECT 74.265 67.620 74.955 67.790 ;
        RECT 73.925 67.000 74.095 67.500 ;
        RECT 75.125 67.000 75.295 67.500 ;
        RECT 74.265 66.710 74.955 66.880 ;
        RECT 74.265 66.120 74.955 66.290 ;
        RECT 73.925 65.500 74.095 66.000 ;
        RECT 75.125 65.500 75.295 66.000 ;
        RECT 74.265 65.210 74.955 65.380 ;
        RECT 75.590 64.720 75.760 78.830 ;
        RECT 73.460 64.550 75.760 64.720 ;
        RECT 76.640 78.680 79.290 78.850 ;
        RECT 76.640 64.820 76.810 78.680 ;
        RECT 77.445 78.120 78.485 78.290 ;
        RECT 77.060 77.500 77.230 78.000 ;
        RECT 78.700 77.500 78.870 78.000 ;
        RECT 77.445 77.210 78.485 77.380 ;
        RECT 77.445 76.620 78.485 76.790 ;
        RECT 77.060 76.000 77.230 76.500 ;
        RECT 78.700 76.000 78.870 76.500 ;
        RECT 77.445 75.710 78.485 75.880 ;
        RECT 77.445 75.120 78.485 75.290 ;
        RECT 77.060 74.500 77.230 75.000 ;
        RECT 78.700 74.500 78.870 75.000 ;
        RECT 77.445 74.210 78.485 74.380 ;
        RECT 77.445 73.620 78.485 73.790 ;
        RECT 77.060 73.000 77.230 73.500 ;
        RECT 78.700 73.000 78.870 73.500 ;
        RECT 77.445 72.710 78.485 72.880 ;
        RECT 77.445 72.120 78.485 72.290 ;
        RECT 77.060 71.500 77.230 72.000 ;
        RECT 78.700 71.500 78.870 72.000 ;
        RECT 77.445 71.210 78.485 71.380 ;
        RECT 77.445 70.620 78.485 70.790 ;
        RECT 77.060 70.000 77.230 70.500 ;
        RECT 78.700 70.000 78.870 70.500 ;
        RECT 77.445 69.710 78.485 69.880 ;
        RECT 77.445 69.120 78.485 69.290 ;
        RECT 77.060 68.500 77.230 69.000 ;
        RECT 78.700 68.500 78.870 69.000 ;
        RECT 77.445 68.210 78.485 68.380 ;
        RECT 77.445 67.620 78.485 67.790 ;
        RECT 77.060 67.000 77.230 67.500 ;
        RECT 78.700 67.000 78.870 67.500 ;
        RECT 77.445 66.710 78.485 66.880 ;
        RECT 77.445 66.120 78.485 66.290 ;
        RECT 77.060 65.500 77.230 66.000 ;
        RECT 78.700 65.500 78.870 66.000 ;
        RECT 77.445 65.210 78.485 65.380 ;
        RECT 79.120 64.820 79.290 78.680 ;
        RECT 76.640 64.650 79.290 64.820 ;
        RECT 80.170 78.830 82.470 79.000 ;
        RECT 80.170 64.720 80.340 78.830 ;
        RECT 80.975 78.120 81.665 78.290 ;
        RECT 80.635 77.500 80.805 78.000 ;
        RECT 81.835 77.500 82.005 78.000 ;
        RECT 80.975 77.210 81.665 77.380 ;
        RECT 80.975 76.620 81.665 76.790 ;
        RECT 80.635 76.000 80.805 76.500 ;
        RECT 81.835 76.000 82.005 76.500 ;
        RECT 80.975 75.710 81.665 75.880 ;
        RECT 80.975 75.120 81.665 75.290 ;
        RECT 80.635 74.500 80.805 75.000 ;
        RECT 81.835 74.500 82.005 75.000 ;
        RECT 80.975 74.210 81.665 74.380 ;
        RECT 80.975 73.620 81.665 73.790 ;
        RECT 80.635 73.000 80.805 73.500 ;
        RECT 81.835 73.000 82.005 73.500 ;
        RECT 80.975 72.710 81.665 72.880 ;
        RECT 80.975 72.120 81.665 72.290 ;
        RECT 80.635 71.500 80.805 72.000 ;
        RECT 81.835 71.500 82.005 72.000 ;
        RECT 80.975 71.210 81.665 71.380 ;
        RECT 80.975 70.620 81.665 70.790 ;
        RECT 80.635 70.000 80.805 70.500 ;
        RECT 81.835 70.000 82.005 70.500 ;
        RECT 80.975 69.710 81.665 69.880 ;
        RECT 80.975 69.120 81.665 69.290 ;
        RECT 80.635 68.500 80.805 69.000 ;
        RECT 81.835 68.500 82.005 69.000 ;
        RECT 80.975 68.210 81.665 68.380 ;
        RECT 80.975 67.620 81.665 67.790 ;
        RECT 80.635 67.000 80.805 67.500 ;
        RECT 81.835 67.000 82.005 67.500 ;
        RECT 80.975 66.710 81.665 66.880 ;
        RECT 80.975 66.120 81.665 66.290 ;
        RECT 80.635 65.500 80.805 66.000 ;
        RECT 81.835 65.500 82.005 66.000 ;
        RECT 80.975 65.210 81.665 65.380 ;
        RECT 82.300 64.720 82.470 78.830 ;
        RECT 80.170 64.550 82.470 64.720 ;
        RECT 83.350 78.680 86.000 78.850 ;
        RECT 83.350 64.820 83.520 78.680 ;
        RECT 84.155 78.120 85.195 78.290 ;
        RECT 83.770 77.500 83.940 78.000 ;
        RECT 85.410 77.500 85.580 78.000 ;
        RECT 84.155 77.210 85.195 77.380 ;
        RECT 84.155 76.620 85.195 76.790 ;
        RECT 83.770 76.000 83.940 76.500 ;
        RECT 85.410 76.000 85.580 76.500 ;
        RECT 84.155 75.710 85.195 75.880 ;
        RECT 84.155 75.120 85.195 75.290 ;
        RECT 83.770 74.500 83.940 75.000 ;
        RECT 85.410 74.500 85.580 75.000 ;
        RECT 84.155 74.210 85.195 74.380 ;
        RECT 84.155 73.620 85.195 73.790 ;
        RECT 83.770 73.000 83.940 73.500 ;
        RECT 85.410 73.000 85.580 73.500 ;
        RECT 84.155 72.710 85.195 72.880 ;
        RECT 84.155 72.120 85.195 72.290 ;
        RECT 83.770 71.500 83.940 72.000 ;
        RECT 85.410 71.500 85.580 72.000 ;
        RECT 84.155 71.210 85.195 71.380 ;
        RECT 84.155 70.620 85.195 70.790 ;
        RECT 83.770 70.000 83.940 70.500 ;
        RECT 85.410 70.000 85.580 70.500 ;
        RECT 84.155 69.710 85.195 69.880 ;
        RECT 84.155 69.120 85.195 69.290 ;
        RECT 83.770 68.500 83.940 69.000 ;
        RECT 85.410 68.500 85.580 69.000 ;
        RECT 84.155 68.210 85.195 68.380 ;
        RECT 84.155 67.620 85.195 67.790 ;
        RECT 83.770 67.000 83.940 67.500 ;
        RECT 85.410 67.000 85.580 67.500 ;
        RECT 84.155 66.710 85.195 66.880 ;
        RECT 84.155 66.120 85.195 66.290 ;
        RECT 83.770 65.500 83.940 66.000 ;
        RECT 85.410 65.500 85.580 66.000 ;
        RECT 84.155 65.210 85.195 65.380 ;
        RECT 85.830 64.820 86.000 78.680 ;
        RECT 83.350 64.650 86.000 64.820 ;
        RECT 86.880 78.830 89.180 79.000 ;
        RECT 86.880 64.720 87.050 78.830 ;
        RECT 87.685 78.120 88.375 78.290 ;
        RECT 87.345 77.500 87.515 78.000 ;
        RECT 88.545 77.500 88.715 78.000 ;
        RECT 87.685 77.210 88.375 77.380 ;
        RECT 87.685 76.620 88.375 76.790 ;
        RECT 87.345 76.000 87.515 76.500 ;
        RECT 88.545 76.000 88.715 76.500 ;
        RECT 87.685 75.710 88.375 75.880 ;
        RECT 87.685 75.120 88.375 75.290 ;
        RECT 87.345 74.500 87.515 75.000 ;
        RECT 88.545 74.500 88.715 75.000 ;
        RECT 87.685 74.210 88.375 74.380 ;
        RECT 87.685 73.620 88.375 73.790 ;
        RECT 87.345 73.000 87.515 73.500 ;
        RECT 88.545 73.000 88.715 73.500 ;
        RECT 87.685 72.710 88.375 72.880 ;
        RECT 87.685 72.120 88.375 72.290 ;
        RECT 87.345 71.500 87.515 72.000 ;
        RECT 88.545 71.500 88.715 72.000 ;
        RECT 87.685 71.210 88.375 71.380 ;
        RECT 87.685 70.620 88.375 70.790 ;
        RECT 87.345 70.000 87.515 70.500 ;
        RECT 88.545 70.000 88.715 70.500 ;
        RECT 87.685 69.710 88.375 69.880 ;
        RECT 87.685 69.120 88.375 69.290 ;
        RECT 87.345 68.500 87.515 69.000 ;
        RECT 88.545 68.500 88.715 69.000 ;
        RECT 87.685 68.210 88.375 68.380 ;
        RECT 87.685 67.620 88.375 67.790 ;
        RECT 87.345 67.000 87.515 67.500 ;
        RECT 88.545 67.000 88.715 67.500 ;
        RECT 87.685 66.710 88.375 66.880 ;
        RECT 87.685 66.120 88.375 66.290 ;
        RECT 87.345 65.500 87.515 66.000 ;
        RECT 88.545 65.500 88.715 66.000 ;
        RECT 87.685 65.210 88.375 65.380 ;
        RECT 89.010 64.720 89.180 78.830 ;
        RECT 86.880 64.550 89.180 64.720 ;
        RECT 90.060 78.680 92.710 78.850 ;
        RECT 90.060 64.820 90.230 78.680 ;
        RECT 90.865 78.120 91.905 78.290 ;
        RECT 90.480 77.500 90.650 78.000 ;
        RECT 92.120 77.500 92.290 78.000 ;
        RECT 90.865 77.210 91.905 77.380 ;
        RECT 90.865 76.620 91.905 76.790 ;
        RECT 90.480 76.000 90.650 76.500 ;
        RECT 92.120 76.000 92.290 76.500 ;
        RECT 90.865 75.710 91.905 75.880 ;
        RECT 90.865 75.120 91.905 75.290 ;
        RECT 90.480 74.500 90.650 75.000 ;
        RECT 92.120 74.500 92.290 75.000 ;
        RECT 90.865 74.210 91.905 74.380 ;
        RECT 90.865 73.620 91.905 73.790 ;
        RECT 90.480 73.000 90.650 73.500 ;
        RECT 92.120 73.000 92.290 73.500 ;
        RECT 90.865 72.710 91.905 72.880 ;
        RECT 90.865 72.120 91.905 72.290 ;
        RECT 90.480 71.500 90.650 72.000 ;
        RECT 92.120 71.500 92.290 72.000 ;
        RECT 90.865 71.210 91.905 71.380 ;
        RECT 90.865 70.620 91.905 70.790 ;
        RECT 90.480 70.000 90.650 70.500 ;
        RECT 92.120 70.000 92.290 70.500 ;
        RECT 90.865 69.710 91.905 69.880 ;
        RECT 90.865 69.120 91.905 69.290 ;
        RECT 90.480 68.500 90.650 69.000 ;
        RECT 92.120 68.500 92.290 69.000 ;
        RECT 90.865 68.210 91.905 68.380 ;
        RECT 90.865 67.620 91.905 67.790 ;
        RECT 90.480 67.000 90.650 67.500 ;
        RECT 92.120 67.000 92.290 67.500 ;
        RECT 90.865 66.710 91.905 66.880 ;
        RECT 90.865 66.120 91.905 66.290 ;
        RECT 90.480 65.500 90.650 66.000 ;
        RECT 92.120 65.500 92.290 66.000 ;
        RECT 90.865 65.210 91.905 65.380 ;
        RECT 92.540 64.820 92.710 78.680 ;
        RECT 90.060 64.650 92.710 64.820 ;
        RECT 93.590 78.830 95.890 79.000 ;
        RECT 93.590 64.720 93.760 78.830 ;
        RECT 94.395 78.120 95.085 78.290 ;
        RECT 94.055 77.500 94.225 78.000 ;
        RECT 95.255 77.500 95.425 78.000 ;
        RECT 94.395 77.210 95.085 77.380 ;
        RECT 94.395 76.620 95.085 76.790 ;
        RECT 94.055 76.000 94.225 76.500 ;
        RECT 95.255 76.000 95.425 76.500 ;
        RECT 94.395 75.710 95.085 75.880 ;
        RECT 94.395 75.120 95.085 75.290 ;
        RECT 94.055 74.500 94.225 75.000 ;
        RECT 95.255 74.500 95.425 75.000 ;
        RECT 94.395 74.210 95.085 74.380 ;
        RECT 94.395 73.620 95.085 73.790 ;
        RECT 94.055 73.000 94.225 73.500 ;
        RECT 95.255 73.000 95.425 73.500 ;
        RECT 94.395 72.710 95.085 72.880 ;
        RECT 94.395 72.120 95.085 72.290 ;
        RECT 94.055 71.500 94.225 72.000 ;
        RECT 95.255 71.500 95.425 72.000 ;
        RECT 94.395 71.210 95.085 71.380 ;
        RECT 94.395 70.620 95.085 70.790 ;
        RECT 94.055 70.000 94.225 70.500 ;
        RECT 95.255 70.000 95.425 70.500 ;
        RECT 94.395 69.710 95.085 69.880 ;
        RECT 94.395 69.120 95.085 69.290 ;
        RECT 94.055 68.500 94.225 69.000 ;
        RECT 95.255 68.500 95.425 69.000 ;
        RECT 94.395 68.210 95.085 68.380 ;
        RECT 94.395 67.620 95.085 67.790 ;
        RECT 94.055 67.000 94.225 67.500 ;
        RECT 95.255 67.000 95.425 67.500 ;
        RECT 94.395 66.710 95.085 66.880 ;
        RECT 94.395 66.120 95.085 66.290 ;
        RECT 94.055 65.500 94.225 66.000 ;
        RECT 95.255 65.500 95.425 66.000 ;
        RECT 94.395 65.210 95.085 65.380 ;
        RECT 95.720 64.720 95.890 78.830 ;
        RECT 93.590 64.550 95.890 64.720 ;
        RECT 96.770 78.680 99.420 78.850 ;
        RECT 96.770 64.820 96.940 78.680 ;
        RECT 97.575 78.120 98.615 78.290 ;
        RECT 97.190 77.500 97.360 78.000 ;
        RECT 98.830 77.500 99.000 78.000 ;
        RECT 97.575 77.210 98.615 77.380 ;
        RECT 97.575 76.620 98.615 76.790 ;
        RECT 97.190 76.000 97.360 76.500 ;
        RECT 98.830 76.000 99.000 76.500 ;
        RECT 97.575 75.710 98.615 75.880 ;
        RECT 97.575 75.120 98.615 75.290 ;
        RECT 97.190 74.500 97.360 75.000 ;
        RECT 98.830 74.500 99.000 75.000 ;
        RECT 97.575 74.210 98.615 74.380 ;
        RECT 97.575 73.620 98.615 73.790 ;
        RECT 97.190 73.000 97.360 73.500 ;
        RECT 98.830 73.000 99.000 73.500 ;
        RECT 97.575 72.710 98.615 72.880 ;
        RECT 97.575 72.120 98.615 72.290 ;
        RECT 97.190 71.500 97.360 72.000 ;
        RECT 98.830 71.500 99.000 72.000 ;
        RECT 97.575 71.210 98.615 71.380 ;
        RECT 97.575 70.620 98.615 70.790 ;
        RECT 97.190 70.000 97.360 70.500 ;
        RECT 98.830 70.000 99.000 70.500 ;
        RECT 97.575 69.710 98.615 69.880 ;
        RECT 97.575 69.120 98.615 69.290 ;
        RECT 97.190 68.500 97.360 69.000 ;
        RECT 98.830 68.500 99.000 69.000 ;
        RECT 97.575 68.210 98.615 68.380 ;
        RECT 97.575 67.620 98.615 67.790 ;
        RECT 97.190 67.000 97.360 67.500 ;
        RECT 98.830 67.000 99.000 67.500 ;
        RECT 97.575 66.710 98.615 66.880 ;
        RECT 97.575 66.120 98.615 66.290 ;
        RECT 97.190 65.500 97.360 66.000 ;
        RECT 98.830 65.500 99.000 66.000 ;
        RECT 97.575 65.210 98.615 65.380 ;
        RECT 99.250 64.820 99.420 78.680 ;
        RECT 96.770 64.650 99.420 64.820 ;
        RECT 100.300 78.830 102.600 79.000 ;
        RECT 100.300 64.720 100.470 78.830 ;
        RECT 101.105 78.120 101.795 78.290 ;
        RECT 100.765 77.500 100.935 78.000 ;
        RECT 101.965 77.500 102.135 78.000 ;
        RECT 101.105 77.210 101.795 77.380 ;
        RECT 101.105 76.620 101.795 76.790 ;
        RECT 100.765 76.000 100.935 76.500 ;
        RECT 101.965 76.000 102.135 76.500 ;
        RECT 101.105 75.710 101.795 75.880 ;
        RECT 101.105 75.120 101.795 75.290 ;
        RECT 100.765 74.500 100.935 75.000 ;
        RECT 101.965 74.500 102.135 75.000 ;
        RECT 101.105 74.210 101.795 74.380 ;
        RECT 101.105 73.620 101.795 73.790 ;
        RECT 100.765 73.000 100.935 73.500 ;
        RECT 101.965 73.000 102.135 73.500 ;
        RECT 101.105 72.710 101.795 72.880 ;
        RECT 101.105 72.120 101.795 72.290 ;
        RECT 100.765 71.500 100.935 72.000 ;
        RECT 101.965 71.500 102.135 72.000 ;
        RECT 101.105 71.210 101.795 71.380 ;
        RECT 101.105 70.620 101.795 70.790 ;
        RECT 100.765 70.000 100.935 70.500 ;
        RECT 101.965 70.000 102.135 70.500 ;
        RECT 101.105 69.710 101.795 69.880 ;
        RECT 101.105 69.120 101.795 69.290 ;
        RECT 100.765 68.500 100.935 69.000 ;
        RECT 101.965 68.500 102.135 69.000 ;
        RECT 101.105 68.210 101.795 68.380 ;
        RECT 101.105 67.620 101.795 67.790 ;
        RECT 100.765 67.000 100.935 67.500 ;
        RECT 101.965 67.000 102.135 67.500 ;
        RECT 101.105 66.710 101.795 66.880 ;
        RECT 101.105 66.120 101.795 66.290 ;
        RECT 100.765 65.500 100.935 66.000 ;
        RECT 101.965 65.500 102.135 66.000 ;
        RECT 101.105 65.210 101.795 65.380 ;
        RECT 102.430 64.720 102.600 78.830 ;
        RECT 100.300 64.550 102.600 64.720 ;
        RECT 111.280 61.285 111.450 164.520 ;
        RECT 27.180 61.115 111.450 61.285 ;
      LAYER met1 ;
        RECT 0.000 224.760 1.000 225.760 ;
        RECT 144.360 224.760 145.360 225.760 ;
        RECT 18.350 207.550 18.850 207.580 ;
        RECT 30.830 207.550 31.330 207.580 ;
        RECT 18.350 207.260 31.330 207.550 ;
        RECT 18.350 207.230 18.970 207.260 ;
        RECT 18.800 206.665 18.970 207.230 ;
        RECT 19.110 206.870 19.570 207.100 ;
        RECT 18.770 205.665 19.000 206.665 ;
        RECT 19.255 206.250 19.425 206.870 ;
        RECT 19.710 206.665 19.880 206.685 ;
        RECT 20.300 206.665 20.470 207.260 ;
        RECT 20.610 206.870 21.070 207.100 ;
        RECT 19.680 206.250 19.910 206.665 ;
        RECT 19.255 206.080 19.910 206.250 ;
        RECT 18.800 205.645 18.970 205.665 ;
        RECT 19.255 205.460 19.425 206.080 ;
        RECT 19.680 205.665 19.910 206.080 ;
        RECT 20.270 205.665 20.500 206.665 ;
        RECT 20.755 206.250 20.925 206.870 ;
        RECT 21.210 206.665 21.380 206.685 ;
        RECT 21.800 206.665 21.970 207.260 ;
        RECT 22.110 206.870 22.570 207.100 ;
        RECT 21.180 206.250 21.410 206.665 ;
        RECT 20.755 206.080 21.410 206.250 ;
        RECT 19.710 205.645 19.880 205.665 ;
        RECT 20.300 205.645 20.470 205.665 ;
        RECT 20.755 205.460 20.925 206.080 ;
        RECT 21.180 205.665 21.410 206.080 ;
        RECT 21.770 205.665 22.000 206.665 ;
        RECT 22.255 206.250 22.425 206.870 ;
        RECT 22.710 206.665 22.880 206.685 ;
        RECT 23.300 206.665 23.470 207.260 ;
        RECT 23.610 206.870 24.070 207.100 ;
        RECT 22.680 206.250 22.910 206.665 ;
        RECT 22.255 206.080 22.910 206.250 ;
        RECT 21.210 205.645 21.380 205.665 ;
        RECT 21.800 205.645 21.970 205.665 ;
        RECT 22.255 205.460 22.425 206.080 ;
        RECT 22.680 205.665 22.910 206.080 ;
        RECT 23.270 205.665 23.500 206.665 ;
        RECT 23.755 206.250 23.925 206.870 ;
        RECT 24.210 206.665 24.380 206.685 ;
        RECT 24.800 206.665 24.970 207.260 ;
        RECT 25.110 206.870 25.570 207.100 ;
        RECT 24.180 206.250 24.410 206.665 ;
        RECT 23.755 206.080 24.410 206.250 ;
        RECT 22.710 205.645 22.880 205.665 ;
        RECT 23.300 205.645 23.470 205.665 ;
        RECT 23.755 205.460 23.925 206.080 ;
        RECT 24.180 205.665 24.410 206.080 ;
        RECT 24.770 205.665 25.000 206.665 ;
        RECT 25.255 206.250 25.425 206.870 ;
        RECT 25.710 206.665 25.880 206.685 ;
        RECT 26.300 206.665 26.470 207.260 ;
        RECT 26.610 206.870 27.070 207.100 ;
        RECT 25.680 206.250 25.910 206.665 ;
        RECT 25.255 206.080 25.910 206.250 ;
        RECT 24.210 205.645 24.380 205.665 ;
        RECT 24.800 205.645 24.970 205.665 ;
        RECT 25.255 205.460 25.425 206.080 ;
        RECT 25.680 205.665 25.910 206.080 ;
        RECT 26.270 205.665 26.500 206.665 ;
        RECT 26.755 206.250 26.925 206.870 ;
        RECT 27.210 206.665 27.380 206.685 ;
        RECT 27.800 206.665 27.970 207.260 ;
        RECT 28.110 206.870 28.570 207.100 ;
        RECT 27.180 206.250 27.410 206.665 ;
        RECT 26.755 206.080 27.410 206.250 ;
        RECT 25.710 205.645 25.880 205.665 ;
        RECT 26.300 205.645 26.470 205.665 ;
        RECT 26.755 205.460 26.925 206.080 ;
        RECT 27.180 205.665 27.410 206.080 ;
        RECT 27.770 205.665 28.000 206.665 ;
        RECT 28.255 206.250 28.425 206.870 ;
        RECT 28.710 206.665 28.880 206.685 ;
        RECT 29.300 206.665 29.470 207.260 ;
        RECT 30.830 207.230 31.330 207.260 ;
        RECT 40.430 207.550 40.930 207.580 ;
        RECT 52.910 207.550 53.410 207.580 ;
        RECT 40.430 207.260 53.410 207.550 ;
        RECT 40.430 207.230 41.050 207.260 ;
        RECT 29.610 206.870 30.070 207.100 ;
        RECT 28.680 206.250 28.910 206.665 ;
        RECT 28.255 206.080 28.910 206.250 ;
        RECT 27.210 205.645 27.380 205.665 ;
        RECT 27.800 205.645 27.970 205.665 ;
        RECT 28.255 205.460 28.425 206.080 ;
        RECT 28.680 205.665 28.910 206.080 ;
        RECT 29.270 205.665 29.500 206.665 ;
        RECT 29.755 206.250 29.925 206.870 ;
        RECT 30.210 206.665 30.380 206.685 ;
        RECT 40.880 206.665 41.050 207.230 ;
        RECT 41.190 206.870 41.650 207.100 ;
        RECT 30.180 206.250 30.410 206.665 ;
        RECT 29.755 206.080 30.410 206.250 ;
        RECT 28.710 205.645 28.880 205.665 ;
        RECT 29.300 205.645 29.470 205.665 ;
        RECT 29.755 205.460 29.925 206.080 ;
        RECT 30.180 205.665 30.410 206.080 ;
        RECT 40.850 205.665 41.080 206.665 ;
        RECT 41.335 206.250 41.505 206.870 ;
        RECT 41.790 206.665 41.960 206.685 ;
        RECT 42.380 206.665 42.550 207.260 ;
        RECT 42.690 206.870 43.150 207.100 ;
        RECT 41.760 206.250 41.990 206.665 ;
        RECT 41.335 206.080 41.990 206.250 ;
        RECT 30.210 205.645 30.380 205.665 ;
        RECT 40.880 205.645 41.050 205.665 ;
        RECT 41.335 205.460 41.505 206.080 ;
        RECT 41.760 205.665 41.990 206.080 ;
        RECT 42.350 205.665 42.580 206.665 ;
        RECT 42.835 206.250 43.005 206.870 ;
        RECT 43.290 206.665 43.460 206.685 ;
        RECT 43.880 206.665 44.050 207.260 ;
        RECT 44.190 206.870 44.650 207.100 ;
        RECT 43.260 206.250 43.490 206.665 ;
        RECT 42.835 206.080 43.490 206.250 ;
        RECT 41.790 205.645 41.960 205.665 ;
        RECT 42.380 205.645 42.550 205.665 ;
        RECT 42.835 205.460 43.005 206.080 ;
        RECT 43.260 205.665 43.490 206.080 ;
        RECT 43.850 205.665 44.080 206.665 ;
        RECT 44.335 206.250 44.505 206.870 ;
        RECT 44.790 206.665 44.960 206.685 ;
        RECT 45.380 206.665 45.550 207.260 ;
        RECT 45.690 206.870 46.150 207.100 ;
        RECT 44.760 206.250 44.990 206.665 ;
        RECT 44.335 206.080 44.990 206.250 ;
        RECT 43.290 205.645 43.460 205.665 ;
        RECT 43.880 205.645 44.050 205.665 ;
        RECT 44.335 205.460 44.505 206.080 ;
        RECT 44.760 205.665 44.990 206.080 ;
        RECT 45.350 205.665 45.580 206.665 ;
        RECT 45.835 206.250 46.005 206.870 ;
        RECT 46.290 206.665 46.460 206.685 ;
        RECT 46.880 206.665 47.050 207.260 ;
        RECT 47.190 206.870 47.650 207.100 ;
        RECT 46.260 206.250 46.490 206.665 ;
        RECT 45.835 206.080 46.490 206.250 ;
        RECT 44.790 205.645 44.960 205.665 ;
        RECT 45.380 205.645 45.550 205.665 ;
        RECT 45.835 205.460 46.005 206.080 ;
        RECT 46.260 205.665 46.490 206.080 ;
        RECT 46.850 205.665 47.080 206.665 ;
        RECT 47.335 206.250 47.505 206.870 ;
        RECT 47.790 206.665 47.960 206.685 ;
        RECT 48.380 206.665 48.550 207.260 ;
        RECT 48.690 206.870 49.150 207.100 ;
        RECT 47.760 206.250 47.990 206.665 ;
        RECT 47.335 206.080 47.990 206.250 ;
        RECT 46.290 205.645 46.460 205.665 ;
        RECT 46.880 205.645 47.050 205.665 ;
        RECT 47.335 205.460 47.505 206.080 ;
        RECT 47.760 205.665 47.990 206.080 ;
        RECT 48.350 205.665 48.580 206.665 ;
        RECT 48.835 206.250 49.005 206.870 ;
        RECT 49.290 206.665 49.460 206.685 ;
        RECT 49.880 206.665 50.050 207.260 ;
        RECT 50.190 206.870 50.650 207.100 ;
        RECT 49.260 206.250 49.490 206.665 ;
        RECT 48.835 206.080 49.490 206.250 ;
        RECT 47.790 205.645 47.960 205.665 ;
        RECT 48.380 205.645 48.550 205.665 ;
        RECT 48.835 205.460 49.005 206.080 ;
        RECT 49.260 205.665 49.490 206.080 ;
        RECT 49.850 205.665 50.080 206.665 ;
        RECT 50.335 206.250 50.505 206.870 ;
        RECT 50.790 206.665 50.960 206.685 ;
        RECT 51.380 206.665 51.550 207.260 ;
        RECT 52.910 207.230 53.410 207.260 ;
        RECT 62.510 207.550 63.010 207.580 ;
        RECT 74.990 207.550 75.490 207.580 ;
        RECT 62.510 207.260 75.490 207.550 ;
        RECT 62.510 207.230 63.130 207.260 ;
        RECT 51.690 206.870 52.150 207.100 ;
        RECT 50.760 206.250 50.990 206.665 ;
        RECT 50.335 206.080 50.990 206.250 ;
        RECT 49.290 205.645 49.460 205.665 ;
        RECT 49.880 205.645 50.050 205.665 ;
        RECT 50.335 205.460 50.505 206.080 ;
        RECT 50.760 205.665 50.990 206.080 ;
        RECT 51.350 205.665 51.580 206.665 ;
        RECT 51.835 206.250 52.005 206.870 ;
        RECT 52.290 206.665 52.460 206.685 ;
        RECT 62.960 206.665 63.130 207.230 ;
        RECT 63.270 206.870 63.730 207.100 ;
        RECT 52.260 206.250 52.490 206.665 ;
        RECT 51.835 206.080 52.490 206.250 ;
        RECT 50.790 205.645 50.960 205.665 ;
        RECT 51.380 205.645 51.550 205.665 ;
        RECT 51.835 205.460 52.005 206.080 ;
        RECT 52.260 205.665 52.490 206.080 ;
        RECT 62.930 205.665 63.160 206.665 ;
        RECT 63.415 206.250 63.585 206.870 ;
        RECT 63.870 206.665 64.040 206.685 ;
        RECT 64.460 206.665 64.630 207.260 ;
        RECT 64.770 206.870 65.230 207.100 ;
        RECT 63.840 206.250 64.070 206.665 ;
        RECT 63.415 206.080 64.070 206.250 ;
        RECT 52.290 205.645 52.460 205.665 ;
        RECT 62.960 205.645 63.130 205.665 ;
        RECT 63.415 205.460 63.585 206.080 ;
        RECT 63.840 205.665 64.070 206.080 ;
        RECT 64.430 205.665 64.660 206.665 ;
        RECT 64.915 206.250 65.085 206.870 ;
        RECT 65.370 206.665 65.540 206.685 ;
        RECT 65.960 206.665 66.130 207.260 ;
        RECT 66.270 206.870 66.730 207.100 ;
        RECT 65.340 206.250 65.570 206.665 ;
        RECT 64.915 206.080 65.570 206.250 ;
        RECT 63.870 205.645 64.040 205.665 ;
        RECT 64.460 205.645 64.630 205.665 ;
        RECT 64.915 205.460 65.085 206.080 ;
        RECT 65.340 205.665 65.570 206.080 ;
        RECT 65.930 205.665 66.160 206.665 ;
        RECT 66.415 206.250 66.585 206.870 ;
        RECT 66.870 206.665 67.040 206.685 ;
        RECT 67.460 206.665 67.630 207.260 ;
        RECT 67.770 206.870 68.230 207.100 ;
        RECT 66.840 206.250 67.070 206.665 ;
        RECT 66.415 206.080 67.070 206.250 ;
        RECT 65.370 205.645 65.540 205.665 ;
        RECT 65.960 205.645 66.130 205.665 ;
        RECT 66.415 205.460 66.585 206.080 ;
        RECT 66.840 205.665 67.070 206.080 ;
        RECT 67.430 205.665 67.660 206.665 ;
        RECT 67.915 206.250 68.085 206.870 ;
        RECT 68.370 206.665 68.540 206.685 ;
        RECT 68.960 206.665 69.130 207.260 ;
        RECT 69.270 206.870 69.730 207.100 ;
        RECT 68.340 206.250 68.570 206.665 ;
        RECT 67.915 206.080 68.570 206.250 ;
        RECT 66.870 205.645 67.040 205.665 ;
        RECT 67.460 205.645 67.630 205.665 ;
        RECT 67.915 205.460 68.085 206.080 ;
        RECT 68.340 205.665 68.570 206.080 ;
        RECT 68.930 205.665 69.160 206.665 ;
        RECT 69.415 206.250 69.585 206.870 ;
        RECT 69.870 206.665 70.040 206.685 ;
        RECT 70.460 206.665 70.630 207.260 ;
        RECT 70.770 206.870 71.230 207.100 ;
        RECT 69.840 206.250 70.070 206.665 ;
        RECT 69.415 206.080 70.070 206.250 ;
        RECT 68.370 205.645 68.540 205.665 ;
        RECT 68.960 205.645 69.130 205.665 ;
        RECT 69.415 205.460 69.585 206.080 ;
        RECT 69.840 205.665 70.070 206.080 ;
        RECT 70.430 205.665 70.660 206.665 ;
        RECT 70.915 206.250 71.085 206.870 ;
        RECT 71.370 206.665 71.540 206.685 ;
        RECT 71.960 206.665 72.130 207.260 ;
        RECT 72.270 206.870 72.730 207.100 ;
        RECT 71.340 206.250 71.570 206.665 ;
        RECT 70.915 206.080 71.570 206.250 ;
        RECT 69.870 205.645 70.040 205.665 ;
        RECT 70.460 205.645 70.630 205.665 ;
        RECT 70.915 205.460 71.085 206.080 ;
        RECT 71.340 205.665 71.570 206.080 ;
        RECT 71.930 205.665 72.160 206.665 ;
        RECT 72.415 206.250 72.585 206.870 ;
        RECT 72.870 206.665 73.040 206.685 ;
        RECT 73.460 206.665 73.630 207.260 ;
        RECT 74.990 207.230 75.490 207.260 ;
        RECT 106.370 207.550 106.870 207.580 ;
        RECT 119.445 207.550 119.945 207.580 ;
        RECT 106.370 207.260 119.945 207.550 ;
        RECT 106.370 207.230 106.870 207.260 ;
        RECT 73.770 206.870 74.230 207.100 ;
        RECT 72.840 206.250 73.070 206.665 ;
        RECT 72.415 206.080 73.070 206.250 ;
        RECT 71.370 205.645 71.540 205.665 ;
        RECT 71.960 205.645 72.130 205.665 ;
        RECT 72.415 205.460 72.585 206.080 ;
        RECT 72.840 205.665 73.070 206.080 ;
        RECT 73.430 205.665 73.660 206.665 ;
        RECT 73.915 206.250 74.085 206.870 ;
        RECT 74.370 206.665 74.540 206.685 ;
        RECT 107.335 206.665 107.505 207.260 ;
        RECT 107.745 207.100 108.005 207.120 ;
        RECT 107.645 206.870 108.105 207.100 ;
        RECT 107.745 206.800 108.005 206.870 ;
        RECT 74.340 206.250 74.570 206.665 ;
        RECT 73.915 206.080 74.570 206.250 ;
        RECT 72.870 205.645 73.040 205.665 ;
        RECT 73.460 205.645 73.630 205.665 ;
        RECT 73.915 205.460 74.085 206.080 ;
        RECT 74.340 205.665 74.570 206.080 ;
        RECT 107.305 205.665 107.535 206.665 ;
        RECT 74.370 205.645 74.540 205.665 ;
        RECT 107.335 205.645 107.505 205.665 ;
        RECT 107.790 205.460 107.960 206.800 ;
        RECT 108.245 206.665 108.415 206.685 ;
        RECT 108.835 206.665 109.005 207.260 ;
        RECT 109.245 207.100 109.505 207.120 ;
        RECT 109.145 206.870 109.605 207.100 ;
        RECT 109.245 206.800 109.505 206.870 ;
        RECT 108.215 205.665 108.445 206.665 ;
        RECT 108.805 205.665 109.035 206.665 ;
        RECT 19.110 205.230 19.570 205.460 ;
        RECT 20.610 205.230 21.070 205.460 ;
        RECT 22.110 205.230 22.570 205.460 ;
        RECT 23.610 205.230 24.070 205.460 ;
        RECT 25.110 205.230 25.570 205.460 ;
        RECT 26.610 205.230 27.070 205.460 ;
        RECT 28.110 205.230 28.570 205.460 ;
        RECT 29.610 205.230 30.070 205.460 ;
        RECT 41.190 205.230 41.650 205.460 ;
        RECT 42.690 205.230 43.150 205.460 ;
        RECT 44.190 205.230 44.650 205.460 ;
        RECT 45.690 205.230 46.150 205.460 ;
        RECT 47.190 205.230 47.650 205.460 ;
        RECT 48.690 205.230 49.150 205.460 ;
        RECT 50.190 205.230 50.650 205.460 ;
        RECT 51.690 205.230 52.150 205.460 ;
        RECT 63.270 205.230 63.730 205.460 ;
        RECT 64.770 205.230 65.230 205.460 ;
        RECT 66.270 205.230 66.730 205.460 ;
        RECT 67.770 205.230 68.230 205.460 ;
        RECT 69.270 205.230 69.730 205.460 ;
        RECT 70.770 205.230 71.230 205.460 ;
        RECT 72.270 205.230 72.730 205.460 ;
        RECT 73.770 205.230 74.230 205.460 ;
        RECT 107.645 205.230 108.105 205.460 ;
        RECT 18.350 204.750 18.850 205.100 ;
        RECT 17.600 203.700 18.850 204.050 ;
        RECT 19.255 203.525 19.425 205.230 ;
        RECT 20.755 203.525 20.925 205.230 ;
        RECT 22.255 203.525 22.425 205.230 ;
        RECT 23.755 203.525 23.925 205.230 ;
        RECT 25.255 203.525 25.425 205.230 ;
        RECT 26.755 203.525 26.925 205.230 ;
        RECT 28.255 203.525 28.425 205.230 ;
        RECT 29.755 203.525 29.925 205.230 ;
        RECT 30.770 204.750 31.330 205.100 ;
        RECT 40.430 204.750 40.930 205.100 ;
        RECT 30.830 203.700 32.080 204.050 ;
        RECT 39.680 203.700 40.930 204.050 ;
        RECT 41.335 203.525 41.505 205.230 ;
        RECT 42.835 203.525 43.005 205.230 ;
        RECT 44.335 203.525 44.505 205.230 ;
        RECT 45.835 203.525 46.005 205.230 ;
        RECT 47.335 203.525 47.505 205.230 ;
        RECT 48.835 203.525 49.005 205.230 ;
        RECT 50.335 203.525 50.505 205.230 ;
        RECT 51.835 203.525 52.005 205.230 ;
        RECT 52.850 204.750 53.410 205.100 ;
        RECT 62.510 204.750 63.010 205.100 ;
        RECT 52.910 203.700 54.160 204.050 ;
        RECT 61.760 203.700 63.010 204.050 ;
        RECT 63.415 203.525 63.585 205.230 ;
        RECT 64.915 203.525 65.085 205.230 ;
        RECT 66.415 203.525 66.585 205.230 ;
        RECT 67.915 203.525 68.085 205.230 ;
        RECT 69.415 203.525 69.585 205.230 ;
        RECT 70.915 203.525 71.085 205.230 ;
        RECT 72.415 203.525 72.585 205.230 ;
        RECT 73.915 203.525 74.085 205.230 ;
        RECT 74.930 204.750 75.490 205.100 ;
        RECT 106.370 204.750 106.870 205.100 ;
        RECT 74.990 203.700 76.240 204.050 ;
        RECT 105.620 203.700 106.870 204.050 ;
        RECT 107.790 203.525 107.960 205.230 ;
        RECT 19.110 203.295 19.570 203.525 ;
        RECT 20.610 203.295 21.070 203.525 ;
        RECT 22.110 203.295 22.570 203.525 ;
        RECT 23.610 203.295 24.070 203.525 ;
        RECT 25.110 203.295 25.570 203.525 ;
        RECT 26.610 203.295 27.070 203.525 ;
        RECT 28.110 203.295 28.570 203.525 ;
        RECT 29.610 203.295 30.070 203.525 ;
        RECT 41.190 203.295 41.650 203.525 ;
        RECT 42.690 203.295 43.150 203.525 ;
        RECT 44.190 203.295 44.650 203.525 ;
        RECT 45.690 203.295 46.150 203.525 ;
        RECT 47.190 203.295 47.650 203.525 ;
        RECT 48.690 203.295 49.150 203.525 ;
        RECT 50.190 203.295 50.650 203.525 ;
        RECT 51.690 203.295 52.150 203.525 ;
        RECT 63.270 203.295 63.730 203.525 ;
        RECT 64.770 203.295 65.230 203.525 ;
        RECT 66.270 203.295 66.730 203.525 ;
        RECT 67.770 203.295 68.230 203.525 ;
        RECT 69.270 203.295 69.730 203.525 ;
        RECT 70.770 203.295 71.230 203.525 ;
        RECT 72.270 203.295 72.730 203.525 ;
        RECT 73.770 203.295 74.230 203.525 ;
        RECT 107.645 203.295 108.105 203.525 ;
        RECT 18.800 203.135 18.970 203.155 ;
        RECT 18.770 202.485 19.000 203.135 ;
        RECT 17.600 201.890 18.100 201.920 ;
        RECT 18.800 201.890 18.970 202.485 ;
        RECT 19.255 202.325 19.425 203.295 ;
        RECT 19.665 202.860 19.925 203.180 ;
        RECT 20.300 203.135 20.470 203.155 ;
        RECT 19.680 202.485 19.910 202.860 ;
        RECT 20.270 202.485 20.500 203.135 ;
        RECT 19.710 202.465 19.880 202.485 ;
        RECT 19.110 202.095 19.570 202.325 ;
        RECT 20.300 201.890 20.470 202.485 ;
        RECT 20.755 202.325 20.925 203.295 ;
        RECT 21.165 202.860 21.425 203.180 ;
        RECT 21.800 203.135 21.970 203.155 ;
        RECT 21.180 202.485 21.410 202.860 ;
        RECT 21.770 202.485 22.000 203.135 ;
        RECT 21.210 202.465 21.380 202.485 ;
        RECT 20.610 202.095 21.070 202.325 ;
        RECT 21.800 201.890 21.970 202.485 ;
        RECT 22.255 202.325 22.425 203.295 ;
        RECT 22.665 202.860 22.925 203.180 ;
        RECT 23.300 203.135 23.470 203.155 ;
        RECT 22.680 202.485 22.910 202.860 ;
        RECT 23.270 202.485 23.500 203.135 ;
        RECT 22.710 202.465 22.880 202.485 ;
        RECT 22.110 202.095 22.570 202.325 ;
        RECT 23.300 201.890 23.470 202.485 ;
        RECT 23.755 202.325 23.925 203.295 ;
        RECT 24.165 202.860 24.425 203.180 ;
        RECT 24.800 203.135 24.970 203.155 ;
        RECT 24.180 202.485 24.410 202.860 ;
        RECT 24.770 202.485 25.000 203.135 ;
        RECT 24.210 202.465 24.380 202.485 ;
        RECT 23.610 202.095 24.070 202.325 ;
        RECT 24.800 201.890 24.970 202.485 ;
        RECT 25.255 202.325 25.425 203.295 ;
        RECT 25.665 202.860 25.925 203.180 ;
        RECT 26.300 203.135 26.470 203.155 ;
        RECT 25.680 202.485 25.910 202.860 ;
        RECT 26.270 202.485 26.500 203.135 ;
        RECT 25.710 202.465 25.880 202.485 ;
        RECT 25.110 202.095 25.570 202.325 ;
        RECT 26.300 201.890 26.470 202.485 ;
        RECT 26.755 202.325 26.925 203.295 ;
        RECT 27.165 202.860 27.425 203.180 ;
        RECT 27.800 203.135 27.970 203.155 ;
        RECT 27.180 202.485 27.410 202.860 ;
        RECT 27.770 202.485 28.000 203.135 ;
        RECT 27.210 202.465 27.380 202.485 ;
        RECT 26.610 202.095 27.070 202.325 ;
        RECT 27.800 201.890 27.970 202.485 ;
        RECT 28.255 202.325 28.425 203.295 ;
        RECT 28.665 202.860 28.925 203.180 ;
        RECT 29.300 203.135 29.470 203.155 ;
        RECT 28.680 202.485 28.910 202.860 ;
        RECT 29.270 202.485 29.500 203.135 ;
        RECT 28.710 202.465 28.880 202.485 ;
        RECT 28.110 202.095 28.570 202.325 ;
        RECT 29.300 201.890 29.470 202.485 ;
        RECT 29.755 202.325 29.925 203.295 ;
        RECT 30.165 202.860 30.425 203.180 ;
        RECT 40.880 203.135 41.050 203.155 ;
        RECT 30.180 202.485 30.410 202.860 ;
        RECT 40.850 202.485 41.080 203.135 ;
        RECT 30.210 202.465 30.380 202.485 ;
        RECT 29.610 202.095 30.070 202.325 ;
        RECT 31.580 201.890 32.080 201.920 ;
        RECT 17.600 201.600 32.080 201.890 ;
        RECT 17.600 201.570 18.100 201.600 ;
        RECT 31.580 201.570 32.080 201.600 ;
        RECT 39.680 201.890 40.180 201.920 ;
        RECT 40.880 201.890 41.050 202.485 ;
        RECT 41.335 202.325 41.505 203.295 ;
        RECT 41.745 202.860 42.005 203.180 ;
        RECT 42.380 203.135 42.550 203.155 ;
        RECT 41.760 202.485 41.990 202.860 ;
        RECT 42.350 202.485 42.580 203.135 ;
        RECT 41.790 202.465 41.960 202.485 ;
        RECT 41.190 202.095 41.650 202.325 ;
        RECT 42.380 201.890 42.550 202.485 ;
        RECT 42.835 202.325 43.005 203.295 ;
        RECT 43.245 202.860 43.505 203.180 ;
        RECT 43.880 203.135 44.050 203.155 ;
        RECT 43.260 202.485 43.490 202.860 ;
        RECT 43.850 202.485 44.080 203.135 ;
        RECT 43.290 202.465 43.460 202.485 ;
        RECT 42.690 202.095 43.150 202.325 ;
        RECT 43.880 201.890 44.050 202.485 ;
        RECT 44.335 202.325 44.505 203.295 ;
        RECT 44.745 202.860 45.005 203.180 ;
        RECT 45.380 203.135 45.550 203.155 ;
        RECT 44.760 202.485 44.990 202.860 ;
        RECT 45.350 202.485 45.580 203.135 ;
        RECT 44.790 202.465 44.960 202.485 ;
        RECT 44.190 202.095 44.650 202.325 ;
        RECT 45.380 201.890 45.550 202.485 ;
        RECT 45.835 202.325 46.005 203.295 ;
        RECT 46.245 202.860 46.505 203.180 ;
        RECT 46.880 203.135 47.050 203.155 ;
        RECT 46.260 202.485 46.490 202.860 ;
        RECT 46.850 202.485 47.080 203.135 ;
        RECT 46.290 202.465 46.460 202.485 ;
        RECT 45.690 202.095 46.150 202.325 ;
        RECT 46.880 201.890 47.050 202.485 ;
        RECT 47.335 202.325 47.505 203.295 ;
        RECT 47.745 202.860 48.005 203.180 ;
        RECT 48.380 203.135 48.550 203.155 ;
        RECT 47.760 202.485 47.990 202.860 ;
        RECT 48.350 202.485 48.580 203.135 ;
        RECT 47.790 202.465 47.960 202.485 ;
        RECT 47.190 202.095 47.650 202.325 ;
        RECT 48.380 201.890 48.550 202.485 ;
        RECT 48.835 202.325 49.005 203.295 ;
        RECT 49.245 202.860 49.505 203.180 ;
        RECT 49.880 203.135 50.050 203.155 ;
        RECT 49.260 202.485 49.490 202.860 ;
        RECT 49.850 202.485 50.080 203.135 ;
        RECT 49.290 202.465 49.460 202.485 ;
        RECT 48.690 202.095 49.150 202.325 ;
        RECT 49.880 201.890 50.050 202.485 ;
        RECT 50.335 202.325 50.505 203.295 ;
        RECT 50.745 202.860 51.005 203.180 ;
        RECT 51.380 203.135 51.550 203.155 ;
        RECT 50.760 202.485 50.990 202.860 ;
        RECT 51.350 202.485 51.580 203.135 ;
        RECT 50.790 202.465 50.960 202.485 ;
        RECT 50.190 202.095 50.650 202.325 ;
        RECT 51.380 201.890 51.550 202.485 ;
        RECT 51.835 202.325 52.005 203.295 ;
        RECT 52.245 202.860 52.505 203.180 ;
        RECT 62.960 203.135 63.130 203.155 ;
        RECT 52.260 202.485 52.490 202.860 ;
        RECT 62.930 202.485 63.160 203.135 ;
        RECT 52.290 202.465 52.460 202.485 ;
        RECT 51.690 202.095 52.150 202.325 ;
        RECT 53.660 201.890 54.160 201.920 ;
        RECT 39.680 201.600 54.160 201.890 ;
        RECT 39.680 201.570 40.180 201.600 ;
        RECT 53.660 201.570 54.160 201.600 ;
        RECT 61.760 201.890 62.260 201.920 ;
        RECT 62.960 201.890 63.130 202.485 ;
        RECT 63.415 202.325 63.585 203.295 ;
        RECT 63.825 202.860 64.085 203.180 ;
        RECT 64.460 203.135 64.630 203.155 ;
        RECT 63.840 202.485 64.070 202.860 ;
        RECT 64.430 202.485 64.660 203.135 ;
        RECT 63.870 202.465 64.040 202.485 ;
        RECT 63.270 202.095 63.730 202.325 ;
        RECT 64.460 201.890 64.630 202.485 ;
        RECT 64.915 202.325 65.085 203.295 ;
        RECT 65.325 202.860 65.585 203.180 ;
        RECT 65.960 203.135 66.130 203.155 ;
        RECT 65.340 202.485 65.570 202.860 ;
        RECT 65.930 202.485 66.160 203.135 ;
        RECT 65.370 202.465 65.540 202.485 ;
        RECT 64.770 202.095 65.230 202.325 ;
        RECT 65.960 201.890 66.130 202.485 ;
        RECT 66.415 202.325 66.585 203.295 ;
        RECT 66.825 202.860 67.085 203.180 ;
        RECT 67.460 203.135 67.630 203.155 ;
        RECT 66.840 202.485 67.070 202.860 ;
        RECT 67.430 202.485 67.660 203.135 ;
        RECT 66.870 202.465 67.040 202.485 ;
        RECT 66.270 202.095 66.730 202.325 ;
        RECT 67.460 201.890 67.630 202.485 ;
        RECT 67.915 202.325 68.085 203.295 ;
        RECT 68.325 202.860 68.585 203.180 ;
        RECT 68.960 203.135 69.130 203.155 ;
        RECT 68.340 202.485 68.570 202.860 ;
        RECT 68.930 202.485 69.160 203.135 ;
        RECT 68.370 202.465 68.540 202.485 ;
        RECT 67.770 202.095 68.230 202.325 ;
        RECT 68.960 201.890 69.130 202.485 ;
        RECT 69.415 202.325 69.585 203.295 ;
        RECT 69.825 202.860 70.085 203.180 ;
        RECT 70.460 203.135 70.630 203.155 ;
        RECT 69.840 202.485 70.070 202.860 ;
        RECT 70.430 202.485 70.660 203.135 ;
        RECT 69.870 202.465 70.040 202.485 ;
        RECT 69.270 202.095 69.730 202.325 ;
        RECT 70.460 201.890 70.630 202.485 ;
        RECT 70.915 202.325 71.085 203.295 ;
        RECT 71.325 202.860 71.585 203.180 ;
        RECT 71.960 203.135 72.130 203.155 ;
        RECT 71.340 202.485 71.570 202.860 ;
        RECT 71.930 202.485 72.160 203.135 ;
        RECT 71.370 202.465 71.540 202.485 ;
        RECT 70.770 202.095 71.230 202.325 ;
        RECT 71.960 201.890 72.130 202.485 ;
        RECT 72.415 202.325 72.585 203.295 ;
        RECT 72.825 202.860 73.085 203.180 ;
        RECT 73.460 203.135 73.630 203.155 ;
        RECT 72.840 202.485 73.070 202.860 ;
        RECT 73.430 202.485 73.660 203.135 ;
        RECT 72.870 202.465 73.040 202.485 ;
        RECT 72.270 202.095 72.730 202.325 ;
        RECT 73.460 201.890 73.630 202.485 ;
        RECT 73.915 202.325 74.085 203.295 ;
        RECT 74.325 202.860 74.585 203.180 ;
        RECT 107.335 203.135 107.505 203.155 ;
        RECT 74.340 202.485 74.570 202.860 ;
        RECT 107.305 202.485 107.535 203.135 ;
        RECT 74.370 202.465 74.540 202.485 ;
        RECT 73.770 202.095 74.230 202.325 ;
        RECT 75.740 201.890 76.240 201.920 ;
        RECT 61.760 201.600 76.240 201.890 ;
        RECT 61.760 201.570 62.260 201.600 ;
        RECT 75.740 201.570 76.240 201.600 ;
        RECT 105.620 201.890 106.120 201.920 ;
        RECT 107.335 201.890 107.505 202.485 ;
        RECT 107.790 202.340 107.960 203.295 ;
        RECT 108.245 203.135 108.415 205.665 ;
        RECT 108.835 205.645 109.005 205.665 ;
        RECT 109.290 205.460 109.460 206.800 ;
        RECT 109.745 206.665 109.915 206.685 ;
        RECT 110.335 206.665 110.505 207.260 ;
        RECT 110.745 207.100 111.005 207.120 ;
        RECT 110.645 206.870 111.105 207.100 ;
        RECT 110.745 206.800 111.005 206.870 ;
        RECT 109.715 205.665 109.945 206.665 ;
        RECT 110.305 205.665 110.535 206.665 ;
        RECT 109.145 205.230 109.605 205.460 ;
        RECT 109.290 203.525 109.460 205.230 ;
        RECT 109.145 203.295 109.605 203.525 ;
        RECT 108.835 203.135 109.005 203.155 ;
        RECT 108.215 202.760 108.445 203.135 ;
        RECT 108.170 202.500 108.490 202.760 ;
        RECT 108.215 202.485 108.445 202.500 ;
        RECT 108.805 202.485 109.035 203.135 ;
        RECT 108.245 202.465 108.415 202.485 ;
        RECT 107.715 202.325 108.035 202.340 ;
        RECT 107.645 202.095 108.105 202.325 ;
        RECT 107.715 202.080 108.035 202.095 ;
        RECT 108.835 201.890 109.005 202.485 ;
        RECT 109.290 202.340 109.460 203.295 ;
        RECT 109.745 203.135 109.915 205.665 ;
        RECT 110.335 205.645 110.505 205.665 ;
        RECT 110.790 205.460 110.960 206.800 ;
        RECT 111.245 206.665 111.415 206.685 ;
        RECT 111.835 206.665 112.005 207.260 ;
        RECT 112.245 207.100 112.505 207.120 ;
        RECT 112.145 206.870 112.605 207.100 ;
        RECT 112.245 206.800 112.505 206.870 ;
        RECT 111.215 205.665 111.445 206.665 ;
        RECT 111.805 205.665 112.035 206.665 ;
        RECT 110.645 205.230 111.105 205.460 ;
        RECT 110.790 203.525 110.960 205.230 ;
        RECT 110.645 203.295 111.105 203.525 ;
        RECT 110.335 203.135 110.505 203.155 ;
        RECT 109.715 202.760 109.945 203.135 ;
        RECT 109.670 202.500 109.990 202.760 ;
        RECT 109.715 202.485 109.945 202.500 ;
        RECT 110.305 202.485 110.535 203.135 ;
        RECT 109.745 202.465 109.915 202.485 ;
        RECT 109.215 202.325 109.535 202.340 ;
        RECT 109.145 202.095 109.605 202.325 ;
        RECT 109.215 202.080 109.535 202.095 ;
        RECT 110.335 201.890 110.505 202.485 ;
        RECT 110.790 202.340 110.960 203.295 ;
        RECT 111.245 203.135 111.415 205.665 ;
        RECT 111.835 205.645 112.005 205.665 ;
        RECT 112.290 205.460 112.460 206.800 ;
        RECT 112.745 206.665 112.915 206.685 ;
        RECT 113.335 206.665 113.505 207.260 ;
        RECT 113.745 207.100 114.005 207.120 ;
        RECT 113.645 206.870 114.105 207.100 ;
        RECT 113.745 206.800 114.005 206.870 ;
        RECT 112.715 205.665 112.945 206.665 ;
        RECT 113.305 205.665 113.535 206.665 ;
        RECT 112.145 205.230 112.605 205.460 ;
        RECT 112.290 203.525 112.460 205.230 ;
        RECT 112.145 203.295 112.605 203.525 ;
        RECT 111.835 203.135 112.005 203.155 ;
        RECT 111.215 202.760 111.445 203.135 ;
        RECT 111.170 202.500 111.490 202.760 ;
        RECT 111.215 202.485 111.445 202.500 ;
        RECT 111.805 202.485 112.035 203.135 ;
        RECT 111.245 202.465 111.415 202.485 ;
        RECT 110.715 202.325 111.035 202.340 ;
        RECT 110.645 202.095 111.105 202.325 ;
        RECT 110.715 202.080 111.035 202.095 ;
        RECT 111.835 201.890 112.005 202.485 ;
        RECT 112.290 202.340 112.460 203.295 ;
        RECT 112.745 203.135 112.915 205.665 ;
        RECT 113.335 205.645 113.505 205.665 ;
        RECT 113.790 205.460 113.960 206.800 ;
        RECT 114.245 206.665 114.415 206.685 ;
        RECT 114.835 206.665 115.005 207.260 ;
        RECT 115.245 207.100 115.505 207.120 ;
        RECT 115.145 206.870 115.605 207.100 ;
        RECT 115.245 206.800 115.505 206.870 ;
        RECT 114.215 205.665 114.445 206.665 ;
        RECT 114.805 205.665 115.035 206.665 ;
        RECT 113.645 205.230 114.105 205.460 ;
        RECT 113.790 203.525 113.960 205.230 ;
        RECT 113.645 203.295 114.105 203.525 ;
        RECT 113.335 203.135 113.505 203.155 ;
        RECT 112.715 202.760 112.945 203.135 ;
        RECT 112.670 202.500 112.990 202.760 ;
        RECT 112.715 202.485 112.945 202.500 ;
        RECT 113.305 202.485 113.535 203.135 ;
        RECT 112.745 202.465 112.915 202.485 ;
        RECT 112.215 202.325 112.535 202.340 ;
        RECT 112.145 202.095 112.605 202.325 ;
        RECT 112.215 202.080 112.535 202.095 ;
        RECT 113.335 201.890 113.505 202.485 ;
        RECT 113.790 202.340 113.960 203.295 ;
        RECT 114.245 203.135 114.415 205.665 ;
        RECT 114.835 205.645 115.005 205.665 ;
        RECT 115.290 205.460 115.460 206.800 ;
        RECT 115.745 206.665 115.915 206.685 ;
        RECT 116.335 206.665 116.505 207.260 ;
        RECT 116.745 207.100 117.005 207.120 ;
        RECT 116.645 206.870 117.105 207.100 ;
        RECT 116.745 206.800 117.005 206.870 ;
        RECT 115.715 205.665 115.945 206.665 ;
        RECT 116.305 205.665 116.535 206.665 ;
        RECT 115.145 205.230 115.605 205.460 ;
        RECT 115.290 203.525 115.460 205.230 ;
        RECT 115.145 203.295 115.605 203.525 ;
        RECT 114.835 203.135 115.005 203.155 ;
        RECT 114.215 202.760 114.445 203.135 ;
        RECT 114.170 202.500 114.490 202.760 ;
        RECT 114.215 202.485 114.445 202.500 ;
        RECT 114.805 202.485 115.035 203.135 ;
        RECT 114.245 202.465 114.415 202.485 ;
        RECT 113.715 202.325 114.035 202.340 ;
        RECT 113.645 202.095 114.105 202.325 ;
        RECT 113.715 202.080 114.035 202.095 ;
        RECT 114.835 201.890 115.005 202.485 ;
        RECT 115.290 202.340 115.460 203.295 ;
        RECT 115.745 203.135 115.915 205.665 ;
        RECT 116.335 205.645 116.505 205.665 ;
        RECT 116.790 205.460 116.960 206.800 ;
        RECT 117.245 206.665 117.415 206.685 ;
        RECT 117.835 206.665 118.005 207.260 ;
        RECT 119.445 207.230 119.945 207.260 ;
        RECT 118.245 207.100 118.505 207.120 ;
        RECT 118.145 206.870 118.605 207.100 ;
        RECT 118.245 206.800 118.505 206.870 ;
        RECT 117.215 205.665 117.445 206.665 ;
        RECT 117.805 205.665 118.035 206.665 ;
        RECT 116.645 205.230 117.105 205.460 ;
        RECT 116.790 203.525 116.960 205.230 ;
        RECT 116.645 203.295 117.105 203.525 ;
        RECT 116.335 203.135 116.505 203.155 ;
        RECT 115.715 202.760 115.945 203.135 ;
        RECT 115.670 202.500 115.990 202.760 ;
        RECT 115.715 202.485 115.945 202.500 ;
        RECT 116.305 202.485 116.535 203.135 ;
        RECT 115.745 202.465 115.915 202.485 ;
        RECT 115.215 202.325 115.535 202.340 ;
        RECT 115.145 202.095 115.605 202.325 ;
        RECT 115.215 202.080 115.535 202.095 ;
        RECT 116.335 201.890 116.505 202.485 ;
        RECT 116.790 202.340 116.960 203.295 ;
        RECT 117.245 203.135 117.415 205.665 ;
        RECT 117.835 205.645 118.005 205.665 ;
        RECT 118.290 205.460 118.460 206.800 ;
        RECT 118.745 206.665 118.915 206.685 ;
        RECT 118.715 205.665 118.945 206.665 ;
        RECT 118.145 205.230 118.605 205.460 ;
        RECT 118.290 203.525 118.460 205.230 ;
        RECT 118.145 203.295 118.605 203.525 ;
        RECT 117.835 203.135 118.005 203.155 ;
        RECT 117.215 202.760 117.445 203.135 ;
        RECT 117.170 202.500 117.490 202.760 ;
        RECT 117.215 202.485 117.445 202.500 ;
        RECT 117.805 202.485 118.035 203.135 ;
        RECT 117.245 202.465 117.415 202.485 ;
        RECT 116.715 202.325 117.035 202.340 ;
        RECT 116.645 202.095 117.105 202.325 ;
        RECT 116.715 202.080 117.035 202.095 ;
        RECT 117.835 201.890 118.005 202.485 ;
        RECT 118.290 202.340 118.460 203.295 ;
        RECT 118.745 203.135 118.915 205.665 ;
        RECT 119.445 204.750 119.945 205.100 ;
        RECT 119.445 203.700 120.695 204.050 ;
        RECT 118.715 202.760 118.945 203.135 ;
        RECT 118.670 202.500 118.990 202.760 ;
        RECT 118.715 202.485 118.945 202.500 ;
        RECT 118.745 202.465 118.915 202.485 ;
        RECT 118.215 202.325 118.535 202.340 ;
        RECT 118.145 202.095 118.605 202.325 ;
        RECT 118.215 202.080 118.535 202.095 ;
        RECT 120.195 201.890 120.695 201.920 ;
        RECT 105.620 201.600 120.695 201.890 ;
        RECT 105.620 201.570 106.120 201.600 ;
        RECT 120.195 201.570 120.695 201.600 ;
        RECT 106.370 200.840 106.870 200.870 ;
        RECT 119.445 200.840 119.945 200.870 ;
        RECT 106.370 200.550 119.945 200.840 ;
        RECT 106.370 200.520 106.870 200.550 ;
        RECT 107.335 199.955 107.505 200.550 ;
        RECT 107.645 200.160 108.105 200.390 ;
        RECT 107.305 198.955 107.535 199.955 ;
        RECT 107.335 198.935 107.505 198.955 ;
        RECT 107.790 198.795 107.960 200.160 ;
        RECT 108.245 199.955 108.415 199.975 ;
        RECT 108.835 199.955 109.005 200.550 ;
        RECT 109.145 200.160 109.605 200.390 ;
        RECT 108.215 198.955 108.445 199.955 ;
        RECT 108.805 198.955 109.035 199.955 ;
        RECT 107.745 198.750 108.005 198.795 ;
        RECT 107.645 198.520 108.105 198.750 ;
        RECT 107.745 198.475 108.005 198.520 ;
        RECT 106.370 198.040 106.870 198.390 ;
        RECT 107.290 197.865 107.550 198.185 ;
        RECT 105.620 196.990 106.870 197.340 ;
        RECT 107.335 196.785 107.505 197.865 ;
        RECT 107.790 197.235 107.960 198.475 ;
        RECT 107.715 196.975 108.035 197.235 ;
        RECT 107.645 196.785 108.105 196.815 ;
        RECT 107.335 196.615 108.105 196.785 ;
        RECT 107.645 196.585 108.105 196.615 ;
        RECT 107.335 196.425 107.505 196.445 ;
        RECT 107.305 195.775 107.535 196.425 ;
        RECT 105.620 195.180 106.120 195.210 ;
        RECT 107.335 195.180 107.505 195.775 ;
        RECT 107.790 195.615 107.960 196.585 ;
        RECT 108.245 196.425 108.415 198.955 ;
        RECT 108.835 198.935 109.005 198.955 ;
        RECT 109.290 198.795 109.460 200.160 ;
        RECT 109.745 199.955 109.915 199.975 ;
        RECT 110.335 199.955 110.505 200.550 ;
        RECT 110.645 200.160 111.105 200.390 ;
        RECT 109.715 198.955 109.945 199.955 ;
        RECT 110.305 198.955 110.535 199.955 ;
        RECT 109.245 198.750 109.505 198.795 ;
        RECT 109.145 198.520 109.605 198.750 ;
        RECT 109.245 198.475 109.505 198.520 ;
        RECT 108.790 197.865 109.050 198.185 ;
        RECT 108.835 196.785 109.005 197.865 ;
        RECT 109.290 197.235 109.460 198.475 ;
        RECT 109.215 196.975 109.535 197.235 ;
        RECT 109.145 196.785 109.605 196.815 ;
        RECT 108.835 196.615 109.605 196.785 ;
        RECT 109.145 196.585 109.605 196.615 ;
        RECT 108.835 196.425 109.005 196.445 ;
        RECT 108.215 196.080 108.445 196.425 ;
        RECT 108.200 195.760 108.460 196.080 ;
        RECT 108.805 195.775 109.035 196.425 ;
        RECT 108.245 195.755 108.415 195.760 ;
        RECT 107.645 195.385 108.105 195.615 ;
        RECT 108.835 195.180 109.005 195.775 ;
        RECT 109.290 195.615 109.460 196.585 ;
        RECT 109.745 196.425 109.915 198.955 ;
        RECT 110.335 198.935 110.505 198.955 ;
        RECT 110.790 198.795 110.960 200.160 ;
        RECT 111.245 199.955 111.415 199.975 ;
        RECT 111.835 199.955 112.005 200.550 ;
        RECT 112.145 200.160 112.605 200.390 ;
        RECT 111.215 198.955 111.445 199.955 ;
        RECT 111.805 198.955 112.035 199.955 ;
        RECT 110.745 198.750 111.005 198.795 ;
        RECT 110.645 198.520 111.105 198.750 ;
        RECT 110.745 198.475 111.005 198.520 ;
        RECT 110.290 197.865 110.550 198.185 ;
        RECT 110.335 196.785 110.505 197.865 ;
        RECT 110.790 197.235 110.960 198.475 ;
        RECT 110.715 196.975 111.035 197.235 ;
        RECT 110.645 196.785 111.105 196.815 ;
        RECT 110.335 196.615 111.105 196.785 ;
        RECT 110.645 196.585 111.105 196.615 ;
        RECT 110.335 196.425 110.505 196.445 ;
        RECT 109.715 196.080 109.945 196.425 ;
        RECT 109.700 195.760 109.960 196.080 ;
        RECT 110.305 195.775 110.535 196.425 ;
        RECT 109.745 195.755 109.915 195.760 ;
        RECT 109.145 195.385 109.605 195.615 ;
        RECT 110.335 195.180 110.505 195.775 ;
        RECT 110.790 195.615 110.960 196.585 ;
        RECT 111.245 196.425 111.415 198.955 ;
        RECT 111.835 198.935 112.005 198.955 ;
        RECT 112.290 198.795 112.460 200.160 ;
        RECT 112.745 199.955 112.915 199.975 ;
        RECT 113.335 199.955 113.505 200.550 ;
        RECT 113.645 200.160 114.105 200.390 ;
        RECT 112.715 198.955 112.945 199.955 ;
        RECT 113.305 198.955 113.535 199.955 ;
        RECT 112.245 198.750 112.505 198.795 ;
        RECT 112.145 198.520 112.605 198.750 ;
        RECT 112.245 198.475 112.505 198.520 ;
        RECT 111.790 197.865 112.050 198.185 ;
        RECT 111.835 196.785 112.005 197.865 ;
        RECT 112.290 197.235 112.460 198.475 ;
        RECT 112.215 196.975 112.535 197.235 ;
        RECT 112.145 196.785 112.605 196.815 ;
        RECT 111.835 196.615 112.605 196.785 ;
        RECT 112.145 196.585 112.605 196.615 ;
        RECT 111.835 196.425 112.005 196.445 ;
        RECT 111.215 196.080 111.445 196.425 ;
        RECT 111.200 195.760 111.460 196.080 ;
        RECT 111.805 195.775 112.035 196.425 ;
        RECT 111.245 195.755 111.415 195.760 ;
        RECT 110.645 195.385 111.105 195.615 ;
        RECT 111.835 195.180 112.005 195.775 ;
        RECT 112.290 195.615 112.460 196.585 ;
        RECT 112.745 196.425 112.915 198.955 ;
        RECT 113.335 198.935 113.505 198.955 ;
        RECT 113.790 198.795 113.960 200.160 ;
        RECT 114.245 199.955 114.415 199.975 ;
        RECT 114.835 199.955 115.005 200.550 ;
        RECT 115.145 200.160 115.605 200.390 ;
        RECT 114.215 198.955 114.445 199.955 ;
        RECT 114.805 198.955 115.035 199.955 ;
        RECT 113.745 198.750 114.005 198.795 ;
        RECT 113.645 198.520 114.105 198.750 ;
        RECT 113.745 198.475 114.005 198.520 ;
        RECT 113.290 197.865 113.550 198.185 ;
        RECT 113.335 196.785 113.505 197.865 ;
        RECT 113.790 197.235 113.960 198.475 ;
        RECT 113.715 196.975 114.035 197.235 ;
        RECT 113.645 196.785 114.105 196.815 ;
        RECT 113.335 196.615 114.105 196.785 ;
        RECT 113.645 196.585 114.105 196.615 ;
        RECT 113.335 196.425 113.505 196.445 ;
        RECT 112.715 196.080 112.945 196.425 ;
        RECT 112.700 195.760 112.960 196.080 ;
        RECT 113.305 195.775 113.535 196.425 ;
        RECT 112.745 195.755 112.915 195.760 ;
        RECT 112.145 195.385 112.605 195.615 ;
        RECT 113.335 195.180 113.505 195.775 ;
        RECT 113.790 195.615 113.960 196.585 ;
        RECT 114.245 196.425 114.415 198.955 ;
        RECT 114.835 198.935 115.005 198.955 ;
        RECT 115.290 198.795 115.460 200.160 ;
        RECT 115.745 199.955 115.915 199.975 ;
        RECT 116.335 199.955 116.505 200.550 ;
        RECT 116.645 200.160 117.105 200.390 ;
        RECT 115.715 198.955 115.945 199.955 ;
        RECT 116.305 198.955 116.535 199.955 ;
        RECT 115.245 198.750 115.505 198.795 ;
        RECT 115.145 198.520 115.605 198.750 ;
        RECT 115.245 198.475 115.505 198.520 ;
        RECT 114.790 197.865 115.050 198.185 ;
        RECT 114.835 196.785 115.005 197.865 ;
        RECT 115.290 197.235 115.460 198.475 ;
        RECT 115.215 196.975 115.535 197.235 ;
        RECT 115.145 196.785 115.605 196.815 ;
        RECT 114.835 196.615 115.605 196.785 ;
        RECT 115.145 196.585 115.605 196.615 ;
        RECT 114.835 196.425 115.005 196.445 ;
        RECT 114.215 196.080 114.445 196.425 ;
        RECT 114.200 195.760 114.460 196.080 ;
        RECT 114.805 195.775 115.035 196.425 ;
        RECT 114.245 195.755 114.415 195.760 ;
        RECT 113.645 195.385 114.105 195.615 ;
        RECT 114.835 195.180 115.005 195.775 ;
        RECT 115.290 195.615 115.460 196.585 ;
        RECT 115.745 196.425 115.915 198.955 ;
        RECT 116.335 198.935 116.505 198.955 ;
        RECT 116.790 198.795 116.960 200.160 ;
        RECT 117.245 199.955 117.415 199.975 ;
        RECT 117.835 199.955 118.005 200.550 ;
        RECT 119.445 200.520 119.945 200.550 ;
        RECT 118.145 200.160 118.605 200.390 ;
        RECT 117.215 198.955 117.445 199.955 ;
        RECT 117.805 198.955 118.035 199.955 ;
        RECT 116.745 198.750 117.005 198.795 ;
        RECT 116.645 198.520 117.105 198.750 ;
        RECT 116.745 198.475 117.005 198.520 ;
        RECT 116.290 197.865 116.550 198.185 ;
        RECT 116.335 196.785 116.505 197.865 ;
        RECT 116.790 197.235 116.960 198.475 ;
        RECT 116.715 196.975 117.035 197.235 ;
        RECT 116.645 196.785 117.105 196.815 ;
        RECT 116.335 196.615 117.105 196.785 ;
        RECT 116.645 196.585 117.105 196.615 ;
        RECT 116.335 196.425 116.505 196.445 ;
        RECT 115.715 196.080 115.945 196.425 ;
        RECT 115.700 195.760 115.960 196.080 ;
        RECT 116.305 195.775 116.535 196.425 ;
        RECT 115.745 195.755 115.915 195.760 ;
        RECT 115.145 195.385 115.605 195.615 ;
        RECT 116.335 195.180 116.505 195.775 ;
        RECT 116.790 195.615 116.960 196.585 ;
        RECT 117.245 196.425 117.415 198.955 ;
        RECT 117.835 198.935 118.005 198.955 ;
        RECT 118.290 198.795 118.460 200.160 ;
        RECT 118.745 199.955 118.915 199.975 ;
        RECT 118.715 198.955 118.945 199.955 ;
        RECT 118.245 198.750 118.505 198.795 ;
        RECT 118.145 198.520 118.605 198.750 ;
        RECT 118.245 198.475 118.505 198.520 ;
        RECT 117.790 197.865 118.050 198.185 ;
        RECT 117.835 196.785 118.005 197.865 ;
        RECT 118.290 197.235 118.460 198.475 ;
        RECT 118.215 196.975 118.535 197.235 ;
        RECT 118.145 196.785 118.605 196.815 ;
        RECT 117.835 196.615 118.605 196.785 ;
        RECT 118.145 196.585 118.605 196.615 ;
        RECT 117.835 196.425 118.005 196.445 ;
        RECT 117.215 196.080 117.445 196.425 ;
        RECT 117.200 195.760 117.460 196.080 ;
        RECT 117.805 195.775 118.035 196.425 ;
        RECT 117.245 195.755 117.415 195.760 ;
        RECT 116.645 195.385 117.105 195.615 ;
        RECT 117.835 195.180 118.005 195.775 ;
        RECT 118.290 195.615 118.460 196.585 ;
        RECT 118.745 196.425 118.915 198.955 ;
        RECT 119.445 198.040 119.945 198.390 ;
        RECT 119.445 196.990 120.695 197.340 ;
        RECT 118.715 196.080 118.945 196.425 ;
        RECT 118.700 195.760 118.960 196.080 ;
        RECT 118.745 195.755 118.915 195.760 ;
        RECT 118.145 195.385 118.605 195.615 ;
        RECT 120.195 195.180 120.695 195.210 ;
        RECT 105.620 194.890 120.695 195.180 ;
        RECT 105.620 194.860 106.120 194.890 ;
        RECT 120.195 194.860 120.695 194.890 ;
        RECT 106.370 194.130 106.870 194.160 ;
        RECT 119.445 194.130 119.945 194.160 ;
        RECT 106.370 193.840 119.945 194.130 ;
        RECT 106.370 193.810 106.870 193.840 ;
        RECT 107.335 193.245 107.505 193.840 ;
        RECT 107.645 193.650 108.105 193.680 ;
        RECT 108.265 193.650 108.585 193.695 ;
        RECT 107.645 193.480 108.585 193.650 ;
        RECT 107.645 193.450 108.105 193.480 ;
        RECT 107.305 192.245 107.535 193.245 ;
        RECT 107.335 192.225 107.505 192.245 ;
        RECT 107.790 192.040 107.960 193.450 ;
        RECT 108.265 193.435 108.585 193.480 ;
        RECT 108.245 193.245 108.415 193.265 ;
        RECT 108.835 193.245 109.005 193.840 ;
        RECT 109.145 193.650 109.605 193.680 ;
        RECT 109.765 193.650 110.085 193.695 ;
        RECT 109.145 193.480 110.085 193.650 ;
        RECT 109.145 193.450 109.605 193.480 ;
        RECT 108.215 193.210 108.445 193.245 ;
        RECT 108.170 192.950 108.490 193.210 ;
        RECT 108.215 192.245 108.445 192.950 ;
        RECT 108.805 192.245 109.035 193.245 ;
        RECT 107.645 191.810 108.105 192.040 ;
        RECT 106.370 191.330 106.870 191.680 ;
        RECT 105.620 190.280 106.870 190.630 ;
        RECT 107.745 190.105 108.005 190.150 ;
        RECT 107.645 189.875 108.105 190.105 ;
        RECT 107.745 189.830 108.005 189.875 ;
        RECT 107.335 189.715 107.505 189.735 ;
        RECT 107.305 189.065 107.535 189.715 ;
        RECT 105.620 188.470 106.120 188.500 ;
        RECT 107.335 188.470 107.505 189.065 ;
        RECT 107.790 188.905 107.960 189.830 ;
        RECT 108.245 189.715 108.415 192.245 ;
        RECT 108.835 192.225 109.005 192.245 ;
        RECT 109.290 192.040 109.460 193.450 ;
        RECT 109.765 193.435 110.085 193.480 ;
        RECT 109.745 193.245 109.915 193.265 ;
        RECT 110.335 193.245 110.505 193.840 ;
        RECT 110.645 193.650 111.105 193.680 ;
        RECT 111.265 193.650 111.585 193.695 ;
        RECT 110.645 193.480 111.585 193.650 ;
        RECT 110.645 193.450 111.105 193.480 ;
        RECT 109.715 193.210 109.945 193.245 ;
        RECT 109.670 192.950 109.990 193.210 ;
        RECT 109.715 192.245 109.945 192.950 ;
        RECT 110.305 192.245 110.535 193.245 ;
        RECT 109.145 191.810 109.605 192.040 ;
        RECT 109.245 190.105 109.505 190.150 ;
        RECT 109.145 189.875 109.605 190.105 ;
        RECT 109.245 189.830 109.505 189.875 ;
        RECT 108.835 189.715 109.005 189.735 ;
        RECT 108.215 189.340 108.445 189.715 ;
        RECT 108.200 189.020 108.460 189.340 ;
        RECT 108.805 189.065 109.035 189.715 ;
        RECT 107.645 188.675 108.105 188.905 ;
        RECT 108.835 188.470 109.005 189.065 ;
        RECT 109.290 188.905 109.460 189.830 ;
        RECT 109.745 189.715 109.915 192.245 ;
        RECT 110.335 192.225 110.505 192.245 ;
        RECT 110.790 192.040 110.960 193.450 ;
        RECT 111.265 193.435 111.585 193.480 ;
        RECT 111.245 193.245 111.415 193.265 ;
        RECT 111.835 193.245 112.005 193.840 ;
        RECT 112.145 193.650 112.605 193.680 ;
        RECT 112.765 193.650 113.085 193.695 ;
        RECT 112.145 193.480 113.085 193.650 ;
        RECT 112.145 193.450 112.605 193.480 ;
        RECT 111.215 193.210 111.445 193.245 ;
        RECT 111.170 192.950 111.490 193.210 ;
        RECT 111.215 192.245 111.445 192.950 ;
        RECT 111.805 192.245 112.035 193.245 ;
        RECT 110.645 191.810 111.105 192.040 ;
        RECT 110.745 190.105 111.005 190.150 ;
        RECT 110.645 189.875 111.105 190.105 ;
        RECT 110.745 189.830 111.005 189.875 ;
        RECT 110.335 189.715 110.505 189.735 ;
        RECT 109.715 189.340 109.945 189.715 ;
        RECT 109.700 189.020 109.960 189.340 ;
        RECT 110.305 189.065 110.535 189.715 ;
        RECT 109.145 188.675 109.605 188.905 ;
        RECT 110.335 188.470 110.505 189.065 ;
        RECT 110.790 188.905 110.960 189.830 ;
        RECT 111.245 189.715 111.415 192.245 ;
        RECT 111.835 192.225 112.005 192.245 ;
        RECT 112.290 192.040 112.460 193.450 ;
        RECT 112.765 193.435 113.085 193.480 ;
        RECT 112.745 193.245 112.915 193.265 ;
        RECT 113.335 193.245 113.505 193.840 ;
        RECT 113.645 193.650 114.105 193.680 ;
        RECT 114.265 193.650 114.585 193.695 ;
        RECT 113.645 193.480 114.585 193.650 ;
        RECT 113.645 193.450 114.105 193.480 ;
        RECT 112.715 193.210 112.945 193.245 ;
        RECT 112.670 192.950 112.990 193.210 ;
        RECT 112.715 192.245 112.945 192.950 ;
        RECT 113.305 192.245 113.535 193.245 ;
        RECT 112.145 191.810 112.605 192.040 ;
        RECT 112.245 190.105 112.505 190.150 ;
        RECT 112.145 189.875 112.605 190.105 ;
        RECT 112.245 189.830 112.505 189.875 ;
        RECT 111.835 189.715 112.005 189.735 ;
        RECT 111.215 189.340 111.445 189.715 ;
        RECT 111.200 189.020 111.460 189.340 ;
        RECT 111.805 189.065 112.035 189.715 ;
        RECT 110.645 188.675 111.105 188.905 ;
        RECT 111.835 188.470 112.005 189.065 ;
        RECT 112.290 188.905 112.460 189.830 ;
        RECT 112.745 189.715 112.915 192.245 ;
        RECT 113.335 192.225 113.505 192.245 ;
        RECT 113.790 192.040 113.960 193.450 ;
        RECT 114.265 193.435 114.585 193.480 ;
        RECT 114.245 193.245 114.415 193.265 ;
        RECT 114.835 193.245 115.005 193.840 ;
        RECT 115.145 193.650 115.605 193.680 ;
        RECT 115.765 193.650 116.085 193.695 ;
        RECT 115.145 193.480 116.085 193.650 ;
        RECT 115.145 193.450 115.605 193.480 ;
        RECT 114.215 193.210 114.445 193.245 ;
        RECT 114.170 192.950 114.490 193.210 ;
        RECT 114.215 192.245 114.445 192.950 ;
        RECT 114.805 192.245 115.035 193.245 ;
        RECT 113.645 191.810 114.105 192.040 ;
        RECT 113.745 190.105 114.005 190.150 ;
        RECT 113.645 189.875 114.105 190.105 ;
        RECT 113.745 189.830 114.005 189.875 ;
        RECT 113.335 189.715 113.505 189.735 ;
        RECT 112.715 189.340 112.945 189.715 ;
        RECT 112.700 189.020 112.960 189.340 ;
        RECT 113.305 189.065 113.535 189.715 ;
        RECT 112.145 188.675 112.605 188.905 ;
        RECT 113.335 188.470 113.505 189.065 ;
        RECT 113.790 188.905 113.960 189.830 ;
        RECT 114.245 189.715 114.415 192.245 ;
        RECT 114.835 192.225 115.005 192.245 ;
        RECT 115.290 192.040 115.460 193.450 ;
        RECT 115.765 193.435 116.085 193.480 ;
        RECT 115.745 193.245 115.915 193.265 ;
        RECT 116.335 193.245 116.505 193.840 ;
        RECT 116.645 193.650 117.105 193.680 ;
        RECT 117.265 193.650 117.585 193.695 ;
        RECT 116.645 193.480 117.585 193.650 ;
        RECT 116.645 193.450 117.105 193.480 ;
        RECT 115.715 193.210 115.945 193.245 ;
        RECT 115.670 192.950 115.990 193.210 ;
        RECT 115.715 192.245 115.945 192.950 ;
        RECT 116.305 192.245 116.535 193.245 ;
        RECT 115.145 191.810 115.605 192.040 ;
        RECT 115.245 190.105 115.505 190.150 ;
        RECT 115.145 189.875 115.605 190.105 ;
        RECT 115.245 189.830 115.505 189.875 ;
        RECT 114.835 189.715 115.005 189.735 ;
        RECT 114.215 189.340 114.445 189.715 ;
        RECT 114.200 189.020 114.460 189.340 ;
        RECT 114.805 189.065 115.035 189.715 ;
        RECT 113.645 188.675 114.105 188.905 ;
        RECT 114.835 188.470 115.005 189.065 ;
        RECT 115.290 188.905 115.460 189.830 ;
        RECT 115.745 189.715 115.915 192.245 ;
        RECT 116.335 192.225 116.505 192.245 ;
        RECT 116.790 192.040 116.960 193.450 ;
        RECT 117.265 193.435 117.585 193.480 ;
        RECT 117.245 193.245 117.415 193.265 ;
        RECT 117.835 193.245 118.005 193.840 ;
        RECT 119.445 193.810 119.945 193.840 ;
        RECT 118.145 193.650 118.605 193.680 ;
        RECT 118.765 193.650 119.085 193.695 ;
        RECT 118.145 193.480 119.085 193.650 ;
        RECT 118.145 193.450 118.605 193.480 ;
        RECT 117.215 193.210 117.445 193.245 ;
        RECT 117.170 192.950 117.490 193.210 ;
        RECT 117.215 192.245 117.445 192.950 ;
        RECT 117.805 192.245 118.035 193.245 ;
        RECT 116.645 191.810 117.105 192.040 ;
        RECT 116.745 190.105 117.005 190.150 ;
        RECT 116.645 189.875 117.105 190.105 ;
        RECT 116.745 189.830 117.005 189.875 ;
        RECT 116.335 189.715 116.505 189.735 ;
        RECT 115.715 189.340 115.945 189.715 ;
        RECT 115.700 189.020 115.960 189.340 ;
        RECT 116.305 189.065 116.535 189.715 ;
        RECT 115.145 188.675 115.605 188.905 ;
        RECT 116.335 188.470 116.505 189.065 ;
        RECT 116.790 188.905 116.960 189.830 ;
        RECT 117.245 189.715 117.415 192.245 ;
        RECT 117.835 192.225 118.005 192.245 ;
        RECT 118.290 192.040 118.460 193.450 ;
        RECT 118.765 193.435 119.085 193.480 ;
        RECT 118.745 193.245 118.915 193.265 ;
        RECT 118.715 193.210 118.945 193.245 ;
        RECT 118.670 192.950 118.990 193.210 ;
        RECT 118.715 192.245 118.945 192.950 ;
        RECT 118.145 191.810 118.605 192.040 ;
        RECT 118.245 190.105 118.505 190.150 ;
        RECT 118.145 189.875 118.605 190.105 ;
        RECT 118.245 189.830 118.505 189.875 ;
        RECT 117.835 189.715 118.005 189.735 ;
        RECT 117.215 189.340 117.445 189.715 ;
        RECT 117.200 189.020 117.460 189.340 ;
        RECT 117.805 189.065 118.035 189.715 ;
        RECT 116.645 188.675 117.105 188.905 ;
        RECT 117.835 188.470 118.005 189.065 ;
        RECT 118.290 188.905 118.460 189.830 ;
        RECT 118.745 189.715 118.915 192.245 ;
        RECT 119.445 191.330 119.945 191.680 ;
        RECT 119.445 190.280 120.695 190.630 ;
        RECT 118.715 189.340 118.945 189.715 ;
        RECT 118.700 189.020 118.960 189.340 ;
        RECT 118.145 188.675 118.605 188.905 ;
        RECT 120.195 188.470 120.695 188.500 ;
        RECT 105.620 188.180 120.695 188.470 ;
        RECT 105.620 188.150 106.120 188.180 ;
        RECT 120.195 188.150 120.695 188.180 ;
        RECT 34.645 163.365 34.945 163.400 ;
        RECT 103.685 163.365 103.985 163.400 ;
        RECT 34.645 163.075 103.985 163.365 ;
        RECT 34.645 163.040 34.945 163.075 ;
        RECT 43.790 162.640 44.250 162.870 ;
        RECT 43.480 162.480 43.650 162.500 ;
        RECT 43.450 161.830 43.680 162.480 ;
        RECT 43.480 160.695 43.650 161.830 ;
        RECT 43.935 161.670 44.105 162.640 ;
        RECT 44.390 162.480 44.560 163.075 ;
        RECT 45.290 162.640 45.750 162.870 ;
        RECT 44.980 162.480 45.150 162.500 ;
        RECT 44.360 161.830 44.590 162.480 ;
        RECT 44.950 161.830 45.180 162.480 ;
        RECT 44.390 161.810 44.560 161.830 ;
        RECT 43.790 161.440 44.250 161.670 ;
        RECT 43.405 160.435 43.725 160.695 ;
        RECT 43.480 159.300 43.650 160.435 ;
        RECT 43.935 160.235 44.105 161.440 ;
        RECT 44.980 160.695 45.150 161.830 ;
        RECT 45.435 161.670 45.605 162.640 ;
        RECT 45.890 162.480 46.060 163.075 ;
        RECT 46.790 162.640 47.250 162.870 ;
        RECT 46.480 162.480 46.650 162.500 ;
        RECT 45.860 161.830 46.090 162.480 ;
        RECT 46.450 161.830 46.680 162.480 ;
        RECT 46.935 162.075 47.105 162.640 ;
        RECT 47.390 162.480 47.560 163.075 ;
        RECT 48.290 162.640 48.750 162.870 ;
        RECT 47.980 162.480 48.150 162.500 ;
        RECT 45.890 161.810 46.060 161.830 ;
        RECT 45.290 161.440 45.750 161.670 ;
        RECT 44.905 160.435 45.225 160.695 ;
        RECT 43.860 159.975 44.180 160.235 ;
        RECT 43.935 159.735 44.105 159.975 ;
        RECT 45.435 159.735 45.605 161.440 ;
        RECT 46.480 160.695 46.650 161.830 ;
        RECT 46.860 161.815 47.180 162.075 ;
        RECT 47.360 161.830 47.590 162.480 ;
        RECT 47.950 161.830 48.180 162.480 ;
        RECT 46.935 161.670 47.105 161.815 ;
        RECT 47.390 161.810 47.560 161.830 ;
        RECT 46.790 161.440 47.250 161.670 ;
        RECT 46.405 160.435 46.725 160.695 ;
        RECT 46.480 160.235 46.650 160.435 ;
        RECT 46.405 159.975 46.725 160.235 ;
        RECT 43.790 159.505 44.250 159.735 ;
        RECT 45.290 159.505 45.750 159.735 ;
        RECT 43.450 158.300 43.680 159.300 ;
        RECT 43.480 158.280 43.650 158.300 ;
        RECT 43.935 158.095 44.105 159.505 ;
        RECT 44.390 159.300 44.560 159.320 ;
        RECT 44.980 159.300 45.150 159.320 ;
        RECT 45.435 159.315 45.605 159.505 ;
        RECT 44.360 158.885 44.590 159.300 ;
        RECT 44.950 158.885 45.180 159.300 ;
        RECT 45.360 159.055 45.680 159.315 ;
        RECT 45.890 159.300 46.060 159.320 ;
        RECT 46.480 159.300 46.650 159.975 ;
        RECT 46.935 159.735 47.105 161.440 ;
        RECT 47.980 160.695 48.150 161.830 ;
        RECT 48.435 161.670 48.605 162.640 ;
        RECT 48.890 162.480 49.060 163.075 ;
        RECT 49.790 162.640 50.250 162.870 ;
        RECT 49.480 162.480 49.650 162.500 ;
        RECT 48.860 161.830 49.090 162.480 ;
        RECT 49.450 161.830 49.680 162.480 ;
        RECT 48.890 161.810 49.060 161.830 ;
        RECT 48.290 161.440 48.750 161.670 ;
        RECT 48.435 161.155 48.605 161.440 ;
        RECT 48.360 160.895 48.680 161.155 ;
        RECT 47.905 160.435 48.225 160.695 ;
        RECT 48.435 159.735 48.605 160.895 ;
        RECT 49.480 160.695 49.650 161.830 ;
        RECT 49.935 161.670 50.105 162.640 ;
        RECT 50.390 162.480 50.560 163.075 ;
        RECT 51.290 162.640 51.750 162.870 ;
        RECT 50.980 162.480 51.150 162.500 ;
        RECT 50.360 161.830 50.590 162.480 ;
        RECT 50.950 161.830 51.180 162.480 ;
        RECT 50.390 161.810 50.560 161.830 ;
        RECT 49.790 161.440 50.250 161.670 ;
        RECT 49.405 160.435 49.725 160.695 ;
        RECT 46.790 159.505 47.250 159.735 ;
        RECT 48.290 159.505 48.750 159.735 ;
        RECT 44.360 158.715 45.180 158.885 ;
        RECT 44.360 158.300 44.590 158.715 ;
        RECT 44.950 158.300 45.180 158.715 ;
        RECT 44.390 158.280 44.560 158.300 ;
        RECT 44.980 158.280 45.150 158.300 ;
        RECT 45.435 158.095 45.605 159.055 ;
        RECT 45.860 158.300 46.090 159.300 ;
        RECT 46.450 158.300 46.680 159.300 ;
        RECT 43.790 157.865 44.250 158.095 ;
        RECT 45.290 157.865 45.750 158.095 ;
        RECT 33.145 157.705 33.445 157.740 ;
        RECT 45.890 157.705 46.060 158.300 ;
        RECT 46.480 158.280 46.650 158.300 ;
        RECT 46.935 158.095 47.105 159.505 ;
        RECT 47.390 159.300 47.560 159.320 ;
        RECT 47.980 159.300 48.150 159.320 ;
        RECT 47.360 158.885 47.590 159.300 ;
        RECT 47.950 158.885 48.180 159.300 ;
        RECT 47.360 158.715 48.180 158.885 ;
        RECT 47.360 158.300 47.590 158.715 ;
        RECT 47.950 158.300 48.180 158.715 ;
        RECT 47.390 158.280 47.560 158.300 ;
        RECT 47.980 158.280 48.150 158.300 ;
        RECT 48.435 158.095 48.605 159.505 ;
        RECT 48.890 159.300 49.060 159.320 ;
        RECT 49.480 159.315 49.650 160.435 ;
        RECT 49.935 160.235 50.105 161.440 ;
        RECT 50.980 160.695 51.150 161.830 ;
        RECT 51.435 161.670 51.605 162.640 ;
        RECT 51.890 162.480 52.060 163.075 ;
        RECT 52.790 162.640 53.250 162.870 ;
        RECT 52.480 162.480 52.650 162.500 ;
        RECT 51.860 161.830 52.090 162.480 ;
        RECT 52.450 162.075 52.680 162.480 ;
        RECT 51.890 161.810 52.060 161.830 ;
        RECT 52.405 161.815 52.725 162.075 ;
        RECT 51.290 161.440 51.750 161.670 ;
        RECT 50.905 160.435 51.225 160.695 ;
        RECT 49.860 159.975 50.180 160.235 ;
        RECT 49.935 159.735 50.105 159.975 ;
        RECT 51.435 159.735 51.605 161.440 ;
        RECT 49.790 159.505 50.250 159.735 ;
        RECT 51.290 159.505 51.750 159.735 ;
        RECT 48.860 158.300 49.090 159.300 ;
        RECT 49.405 159.055 49.725 159.315 ;
        RECT 49.450 158.300 49.680 159.055 ;
        RECT 46.790 157.865 47.250 158.095 ;
        RECT 48.290 157.865 48.750 158.095 ;
        RECT 48.890 157.705 49.060 158.300 ;
        RECT 49.480 158.280 49.650 158.300 ;
        RECT 49.935 158.095 50.105 159.505 ;
        RECT 50.390 159.300 50.560 159.320 ;
        RECT 50.980 159.300 51.150 159.320 ;
        RECT 51.435 159.315 51.605 159.505 ;
        RECT 50.360 158.885 50.590 159.300 ;
        RECT 50.950 158.885 51.180 159.300 ;
        RECT 51.360 159.055 51.680 159.315 ;
        RECT 51.890 159.300 52.060 159.320 ;
        RECT 52.480 159.300 52.650 161.815 ;
        RECT 52.935 161.670 53.105 162.640 ;
        RECT 53.390 162.480 53.560 163.075 ;
        RECT 54.360 162.870 54.680 162.885 ;
        RECT 54.290 162.640 54.750 162.870 ;
        RECT 54.360 162.625 54.680 162.640 ;
        RECT 53.980 162.480 54.150 162.500 ;
        RECT 53.360 161.830 53.590 162.480 ;
        RECT 53.950 161.830 54.180 162.480 ;
        RECT 53.390 161.810 53.560 161.830 ;
        RECT 52.790 161.440 53.250 161.670 ;
        RECT 52.935 160.235 53.105 161.440 ;
        RECT 53.980 161.155 54.150 161.830 ;
        RECT 54.435 161.670 54.605 162.625 ;
        RECT 54.890 162.480 55.060 163.075 ;
        RECT 57.270 162.640 57.730 162.870 ;
        RECT 56.960 162.480 57.130 162.500 ;
        RECT 54.860 161.830 55.090 162.480 ;
        RECT 56.930 161.830 57.160 162.480 ;
        RECT 54.890 161.810 55.060 161.830 ;
        RECT 54.290 161.440 54.750 161.670 ;
        RECT 53.905 160.895 54.225 161.155 ;
        RECT 52.860 159.975 53.180 160.235 ;
        RECT 52.935 159.735 53.105 159.975 ;
        RECT 52.790 159.505 53.250 159.735 ;
        RECT 50.360 158.715 51.180 158.885 ;
        RECT 50.360 158.300 50.590 158.715 ;
        RECT 50.950 158.300 51.180 158.715 ;
        RECT 50.390 158.280 50.560 158.300 ;
        RECT 50.980 158.280 51.150 158.300 ;
        RECT 51.435 158.095 51.605 159.055 ;
        RECT 51.860 158.300 52.090 159.300 ;
        RECT 52.450 158.300 52.680 159.300 ;
        RECT 49.790 157.865 50.250 158.095 ;
        RECT 51.290 157.865 51.750 158.095 ;
        RECT 51.890 157.705 52.060 158.300 ;
        RECT 52.480 158.280 52.650 158.300 ;
        RECT 52.935 158.095 53.105 159.505 ;
        RECT 53.390 159.300 53.560 159.320 ;
        RECT 53.980 159.300 54.150 160.895 ;
        RECT 54.435 159.735 54.605 161.440 ;
        RECT 56.960 160.695 57.130 161.830 ;
        RECT 57.415 161.670 57.585 162.640 ;
        RECT 57.870 162.480 58.040 163.075 ;
        RECT 58.770 162.640 59.230 162.870 ;
        RECT 58.460 162.480 58.630 162.500 ;
        RECT 57.840 161.830 58.070 162.480 ;
        RECT 58.430 161.830 58.660 162.480 ;
        RECT 57.870 161.810 58.040 161.830 ;
        RECT 57.270 161.440 57.730 161.670 ;
        RECT 56.885 160.435 57.205 160.695 ;
        RECT 54.290 159.505 54.750 159.735 ;
        RECT 54.435 159.315 54.605 159.505 ;
        RECT 53.360 158.300 53.590 159.300 ;
        RECT 53.950 158.300 54.180 159.300 ;
        RECT 54.360 159.055 54.680 159.315 ;
        RECT 54.890 159.300 55.060 159.320 ;
        RECT 56.960 159.300 57.130 160.435 ;
        RECT 57.415 160.235 57.585 161.440 ;
        RECT 58.460 160.695 58.630 161.830 ;
        RECT 58.915 161.670 59.085 162.640 ;
        RECT 59.370 162.480 59.540 163.075 ;
        RECT 60.270 162.640 60.730 162.870 ;
        RECT 59.960 162.480 60.130 162.500 ;
        RECT 59.340 161.830 59.570 162.480 ;
        RECT 59.930 161.830 60.160 162.480 ;
        RECT 60.415 162.075 60.585 162.640 ;
        RECT 60.870 162.480 61.040 163.075 ;
        RECT 61.770 162.640 62.230 162.870 ;
        RECT 61.460 162.480 61.630 162.500 ;
        RECT 59.370 161.810 59.540 161.830 ;
        RECT 58.770 161.440 59.230 161.670 ;
        RECT 58.385 160.435 58.705 160.695 ;
        RECT 57.340 159.975 57.660 160.235 ;
        RECT 57.415 159.735 57.585 159.975 ;
        RECT 58.915 159.735 59.085 161.440 ;
        RECT 59.960 160.695 60.130 161.830 ;
        RECT 60.340 161.815 60.660 162.075 ;
        RECT 60.840 161.830 61.070 162.480 ;
        RECT 61.430 161.830 61.660 162.480 ;
        RECT 60.415 161.670 60.585 161.815 ;
        RECT 60.870 161.810 61.040 161.830 ;
        RECT 60.270 161.440 60.730 161.670 ;
        RECT 59.885 160.435 60.205 160.695 ;
        RECT 59.960 160.235 60.130 160.435 ;
        RECT 59.885 159.975 60.205 160.235 ;
        RECT 57.270 159.505 57.730 159.735 ;
        RECT 58.770 159.505 59.230 159.735 ;
        RECT 52.790 157.865 53.250 158.095 ;
        RECT 53.390 157.705 53.560 158.300 ;
        RECT 53.980 158.280 54.150 158.300 ;
        RECT 54.435 158.095 54.605 159.055 ;
        RECT 54.860 158.300 55.090 159.300 ;
        RECT 56.930 158.300 57.160 159.300 ;
        RECT 54.290 157.865 54.750 158.095 ;
        RECT 54.890 157.705 55.060 158.300 ;
        RECT 56.960 158.280 57.130 158.300 ;
        RECT 57.415 158.095 57.585 159.505 ;
        RECT 57.870 159.300 58.040 159.320 ;
        RECT 58.460 159.300 58.630 159.320 ;
        RECT 58.915 159.315 59.085 159.505 ;
        RECT 57.840 158.885 58.070 159.300 ;
        RECT 58.430 158.885 58.660 159.300 ;
        RECT 58.840 159.055 59.160 159.315 ;
        RECT 59.370 159.300 59.540 159.320 ;
        RECT 59.960 159.300 60.130 159.975 ;
        RECT 60.415 159.735 60.585 161.440 ;
        RECT 61.460 160.695 61.630 161.830 ;
        RECT 61.915 161.670 62.085 162.640 ;
        RECT 62.370 162.480 62.540 163.075 ;
        RECT 63.270 162.640 63.730 162.870 ;
        RECT 62.960 162.480 63.130 162.500 ;
        RECT 62.340 161.830 62.570 162.480 ;
        RECT 62.930 161.830 63.160 162.480 ;
        RECT 62.370 161.810 62.540 161.830 ;
        RECT 61.770 161.440 62.230 161.670 ;
        RECT 61.915 161.155 62.085 161.440 ;
        RECT 61.840 160.895 62.160 161.155 ;
        RECT 61.385 160.435 61.705 160.695 ;
        RECT 61.915 159.735 62.085 160.895 ;
        RECT 62.960 160.695 63.130 161.830 ;
        RECT 63.415 161.670 63.585 162.640 ;
        RECT 63.870 162.480 64.040 163.075 ;
        RECT 64.770 162.640 65.230 162.870 ;
        RECT 64.460 162.480 64.630 162.500 ;
        RECT 63.840 161.830 64.070 162.480 ;
        RECT 64.430 161.830 64.660 162.480 ;
        RECT 63.870 161.810 64.040 161.830 ;
        RECT 63.270 161.440 63.730 161.670 ;
        RECT 62.885 160.435 63.205 160.695 ;
        RECT 60.270 159.505 60.730 159.735 ;
        RECT 61.770 159.505 62.230 159.735 ;
        RECT 57.840 158.715 58.660 158.885 ;
        RECT 57.840 158.300 58.070 158.715 ;
        RECT 58.430 158.300 58.660 158.715 ;
        RECT 57.870 158.280 58.040 158.300 ;
        RECT 58.460 158.280 58.630 158.300 ;
        RECT 58.915 158.095 59.085 159.055 ;
        RECT 59.340 158.300 59.570 159.300 ;
        RECT 59.930 158.300 60.160 159.300 ;
        RECT 57.270 157.865 57.730 158.095 ;
        RECT 58.770 157.865 59.230 158.095 ;
        RECT 59.370 157.705 59.540 158.300 ;
        RECT 59.960 158.280 60.130 158.300 ;
        RECT 60.415 158.095 60.585 159.505 ;
        RECT 60.870 159.300 61.040 159.320 ;
        RECT 61.460 159.300 61.630 159.320 ;
        RECT 60.840 158.885 61.070 159.300 ;
        RECT 61.430 158.885 61.660 159.300 ;
        RECT 60.840 158.715 61.660 158.885 ;
        RECT 60.840 158.300 61.070 158.715 ;
        RECT 61.430 158.300 61.660 158.715 ;
        RECT 60.870 158.280 61.040 158.300 ;
        RECT 61.460 158.280 61.630 158.300 ;
        RECT 61.915 158.095 62.085 159.505 ;
        RECT 62.370 159.300 62.540 159.320 ;
        RECT 62.960 159.315 63.130 160.435 ;
        RECT 63.415 160.235 63.585 161.440 ;
        RECT 64.460 160.695 64.630 161.830 ;
        RECT 64.915 161.670 65.085 162.640 ;
        RECT 65.370 162.480 65.540 163.075 ;
        RECT 66.270 162.640 66.730 162.870 ;
        RECT 65.960 162.480 66.130 162.500 ;
        RECT 65.340 161.830 65.570 162.480 ;
        RECT 65.930 162.075 66.160 162.480 ;
        RECT 65.370 161.810 65.540 161.830 ;
        RECT 65.885 161.815 66.205 162.075 ;
        RECT 64.770 161.440 65.230 161.670 ;
        RECT 64.385 160.435 64.705 160.695 ;
        RECT 63.340 159.975 63.660 160.235 ;
        RECT 63.415 159.735 63.585 159.975 ;
        RECT 64.915 159.735 65.085 161.440 ;
        RECT 63.270 159.505 63.730 159.735 ;
        RECT 64.770 159.505 65.230 159.735 ;
        RECT 62.340 158.300 62.570 159.300 ;
        RECT 62.885 159.055 63.205 159.315 ;
        RECT 62.930 158.300 63.160 159.055 ;
        RECT 60.270 157.865 60.730 158.095 ;
        RECT 61.770 157.865 62.230 158.095 ;
        RECT 62.370 157.705 62.540 158.300 ;
        RECT 62.960 158.280 63.130 158.300 ;
        RECT 63.415 158.095 63.585 159.505 ;
        RECT 63.870 159.300 64.040 159.320 ;
        RECT 64.460 159.300 64.630 159.320 ;
        RECT 64.915 159.315 65.085 159.505 ;
        RECT 63.840 158.885 64.070 159.300 ;
        RECT 64.430 158.885 64.660 159.300 ;
        RECT 64.840 159.055 65.160 159.315 ;
        RECT 65.370 159.300 65.540 159.320 ;
        RECT 65.960 159.300 66.130 161.815 ;
        RECT 66.415 161.670 66.585 162.640 ;
        RECT 66.870 162.480 67.040 163.075 ;
        RECT 67.840 162.870 68.160 162.885 ;
        RECT 67.770 162.640 68.230 162.870 ;
        RECT 67.840 162.625 68.160 162.640 ;
        RECT 67.460 162.480 67.630 162.500 ;
        RECT 66.840 161.830 67.070 162.480 ;
        RECT 67.430 161.830 67.660 162.480 ;
        RECT 66.870 161.810 67.040 161.830 ;
        RECT 66.270 161.440 66.730 161.670 ;
        RECT 66.415 160.235 66.585 161.440 ;
        RECT 67.460 161.155 67.630 161.830 ;
        RECT 67.915 161.670 68.085 162.625 ;
        RECT 68.370 162.480 68.540 163.075 ;
        RECT 70.750 162.640 71.210 162.870 ;
        RECT 70.440 162.480 70.610 162.500 ;
        RECT 68.340 161.830 68.570 162.480 ;
        RECT 70.410 161.830 70.640 162.480 ;
        RECT 68.370 161.810 68.540 161.830 ;
        RECT 67.770 161.440 68.230 161.670 ;
        RECT 67.385 160.895 67.705 161.155 ;
        RECT 66.340 159.975 66.660 160.235 ;
        RECT 66.415 159.735 66.585 159.975 ;
        RECT 66.270 159.505 66.730 159.735 ;
        RECT 63.840 158.715 64.660 158.885 ;
        RECT 63.840 158.300 64.070 158.715 ;
        RECT 64.430 158.300 64.660 158.715 ;
        RECT 63.870 158.280 64.040 158.300 ;
        RECT 64.460 158.280 64.630 158.300 ;
        RECT 64.915 158.095 65.085 159.055 ;
        RECT 65.340 158.300 65.570 159.300 ;
        RECT 65.930 158.300 66.160 159.300 ;
        RECT 63.270 157.865 63.730 158.095 ;
        RECT 64.770 157.865 65.230 158.095 ;
        RECT 65.370 157.705 65.540 158.300 ;
        RECT 65.960 158.280 66.130 158.300 ;
        RECT 66.415 158.095 66.585 159.505 ;
        RECT 66.870 159.300 67.040 159.320 ;
        RECT 67.460 159.300 67.630 160.895 ;
        RECT 67.915 159.735 68.085 161.440 ;
        RECT 70.440 160.695 70.610 161.830 ;
        RECT 70.895 161.670 71.065 162.640 ;
        RECT 71.350 162.480 71.520 163.075 ;
        RECT 72.250 162.640 72.710 162.870 ;
        RECT 71.940 162.480 72.110 162.500 ;
        RECT 71.320 161.830 71.550 162.480 ;
        RECT 71.910 161.830 72.140 162.480 ;
        RECT 71.350 161.810 71.520 161.830 ;
        RECT 70.750 161.440 71.210 161.670 ;
        RECT 70.365 160.435 70.685 160.695 ;
        RECT 67.770 159.505 68.230 159.735 ;
        RECT 67.915 159.315 68.085 159.505 ;
        RECT 66.840 158.300 67.070 159.300 ;
        RECT 67.430 158.300 67.660 159.300 ;
        RECT 67.840 159.055 68.160 159.315 ;
        RECT 68.370 159.300 68.540 159.320 ;
        RECT 70.440 159.300 70.610 160.435 ;
        RECT 70.895 160.235 71.065 161.440 ;
        RECT 71.940 160.695 72.110 161.830 ;
        RECT 72.395 161.670 72.565 162.640 ;
        RECT 72.850 162.480 73.020 163.075 ;
        RECT 73.750 162.640 74.210 162.870 ;
        RECT 73.440 162.480 73.610 162.500 ;
        RECT 72.820 161.830 73.050 162.480 ;
        RECT 73.410 161.830 73.640 162.480 ;
        RECT 73.895 162.075 74.065 162.640 ;
        RECT 74.350 162.480 74.520 163.075 ;
        RECT 75.250 162.640 75.710 162.870 ;
        RECT 74.940 162.480 75.110 162.500 ;
        RECT 72.850 161.810 73.020 161.830 ;
        RECT 72.250 161.440 72.710 161.670 ;
        RECT 71.865 160.435 72.185 160.695 ;
        RECT 70.820 159.975 71.140 160.235 ;
        RECT 70.895 159.735 71.065 159.975 ;
        RECT 72.395 159.735 72.565 161.440 ;
        RECT 73.440 160.695 73.610 161.830 ;
        RECT 73.820 161.815 74.140 162.075 ;
        RECT 74.320 161.830 74.550 162.480 ;
        RECT 74.910 161.830 75.140 162.480 ;
        RECT 73.895 161.670 74.065 161.815 ;
        RECT 74.350 161.810 74.520 161.830 ;
        RECT 73.750 161.440 74.210 161.670 ;
        RECT 73.365 160.435 73.685 160.695 ;
        RECT 73.440 160.235 73.610 160.435 ;
        RECT 73.365 159.975 73.685 160.235 ;
        RECT 70.750 159.505 71.210 159.735 ;
        RECT 72.250 159.505 72.710 159.735 ;
        RECT 66.270 157.865 66.730 158.095 ;
        RECT 66.870 157.705 67.040 158.300 ;
        RECT 67.460 158.280 67.630 158.300 ;
        RECT 67.915 158.095 68.085 159.055 ;
        RECT 68.340 158.300 68.570 159.300 ;
        RECT 70.410 158.300 70.640 159.300 ;
        RECT 67.770 157.865 68.230 158.095 ;
        RECT 68.370 157.705 68.540 158.300 ;
        RECT 70.440 158.280 70.610 158.300 ;
        RECT 70.895 158.095 71.065 159.505 ;
        RECT 71.350 159.300 71.520 159.320 ;
        RECT 71.940 159.300 72.110 159.320 ;
        RECT 72.395 159.315 72.565 159.505 ;
        RECT 71.320 158.885 71.550 159.300 ;
        RECT 71.910 158.885 72.140 159.300 ;
        RECT 72.320 159.055 72.640 159.315 ;
        RECT 72.850 159.300 73.020 159.320 ;
        RECT 73.440 159.300 73.610 159.975 ;
        RECT 73.895 159.735 74.065 161.440 ;
        RECT 74.940 160.695 75.110 161.830 ;
        RECT 75.395 161.670 75.565 162.640 ;
        RECT 75.850 162.480 76.020 163.075 ;
        RECT 76.750 162.640 77.210 162.870 ;
        RECT 76.440 162.480 76.610 162.500 ;
        RECT 75.820 161.830 76.050 162.480 ;
        RECT 76.410 161.830 76.640 162.480 ;
        RECT 75.850 161.810 76.020 161.830 ;
        RECT 75.250 161.440 75.710 161.670 ;
        RECT 75.395 161.155 75.565 161.440 ;
        RECT 75.320 160.895 75.640 161.155 ;
        RECT 74.865 160.435 75.185 160.695 ;
        RECT 75.395 159.735 75.565 160.895 ;
        RECT 76.440 160.695 76.610 161.830 ;
        RECT 76.895 161.670 77.065 162.640 ;
        RECT 77.350 162.480 77.520 163.075 ;
        RECT 78.250 162.640 78.710 162.870 ;
        RECT 77.940 162.480 78.110 162.500 ;
        RECT 77.320 161.830 77.550 162.480 ;
        RECT 77.910 161.830 78.140 162.480 ;
        RECT 77.350 161.810 77.520 161.830 ;
        RECT 76.750 161.440 77.210 161.670 ;
        RECT 76.365 160.435 76.685 160.695 ;
        RECT 73.750 159.505 74.210 159.735 ;
        RECT 75.250 159.505 75.710 159.735 ;
        RECT 71.320 158.715 72.140 158.885 ;
        RECT 71.320 158.300 71.550 158.715 ;
        RECT 71.910 158.300 72.140 158.715 ;
        RECT 71.350 158.280 71.520 158.300 ;
        RECT 71.940 158.280 72.110 158.300 ;
        RECT 72.395 158.095 72.565 159.055 ;
        RECT 72.820 158.300 73.050 159.300 ;
        RECT 73.410 158.300 73.640 159.300 ;
        RECT 70.750 157.865 71.210 158.095 ;
        RECT 72.250 157.865 72.710 158.095 ;
        RECT 72.850 157.705 73.020 158.300 ;
        RECT 73.440 158.280 73.610 158.300 ;
        RECT 73.895 158.095 74.065 159.505 ;
        RECT 74.350 159.300 74.520 159.320 ;
        RECT 74.940 159.300 75.110 159.320 ;
        RECT 74.320 158.885 74.550 159.300 ;
        RECT 74.910 158.885 75.140 159.300 ;
        RECT 74.320 158.715 75.140 158.885 ;
        RECT 74.320 158.300 74.550 158.715 ;
        RECT 74.910 158.300 75.140 158.715 ;
        RECT 74.350 158.280 74.520 158.300 ;
        RECT 74.940 158.280 75.110 158.300 ;
        RECT 75.395 158.095 75.565 159.505 ;
        RECT 75.850 159.300 76.020 159.320 ;
        RECT 76.440 159.315 76.610 160.435 ;
        RECT 76.895 160.235 77.065 161.440 ;
        RECT 77.940 160.695 78.110 161.830 ;
        RECT 78.395 161.670 78.565 162.640 ;
        RECT 78.850 162.480 79.020 163.075 ;
        RECT 79.750 162.640 80.210 162.870 ;
        RECT 79.440 162.480 79.610 162.500 ;
        RECT 78.820 161.830 79.050 162.480 ;
        RECT 79.410 162.075 79.640 162.480 ;
        RECT 78.850 161.810 79.020 161.830 ;
        RECT 79.365 161.815 79.685 162.075 ;
        RECT 78.250 161.440 78.710 161.670 ;
        RECT 77.865 160.435 78.185 160.695 ;
        RECT 76.820 159.975 77.140 160.235 ;
        RECT 76.895 159.735 77.065 159.975 ;
        RECT 78.395 159.735 78.565 161.440 ;
        RECT 76.750 159.505 77.210 159.735 ;
        RECT 78.250 159.505 78.710 159.735 ;
        RECT 75.820 158.300 76.050 159.300 ;
        RECT 76.365 159.055 76.685 159.315 ;
        RECT 76.410 158.300 76.640 159.055 ;
        RECT 73.750 157.865 74.210 158.095 ;
        RECT 75.250 157.865 75.710 158.095 ;
        RECT 75.850 157.705 76.020 158.300 ;
        RECT 76.440 158.280 76.610 158.300 ;
        RECT 76.895 158.095 77.065 159.505 ;
        RECT 77.350 159.300 77.520 159.320 ;
        RECT 77.940 159.300 78.110 159.320 ;
        RECT 78.395 159.315 78.565 159.505 ;
        RECT 77.320 158.885 77.550 159.300 ;
        RECT 77.910 158.885 78.140 159.300 ;
        RECT 78.320 159.055 78.640 159.315 ;
        RECT 78.850 159.300 79.020 159.320 ;
        RECT 79.440 159.300 79.610 161.815 ;
        RECT 79.895 161.670 80.065 162.640 ;
        RECT 80.350 162.480 80.520 163.075 ;
        RECT 81.320 162.870 81.640 162.885 ;
        RECT 81.250 162.640 81.710 162.870 ;
        RECT 81.320 162.625 81.640 162.640 ;
        RECT 80.940 162.480 81.110 162.500 ;
        RECT 80.320 161.830 80.550 162.480 ;
        RECT 80.910 161.830 81.140 162.480 ;
        RECT 80.350 161.810 80.520 161.830 ;
        RECT 79.750 161.440 80.210 161.670 ;
        RECT 79.895 160.235 80.065 161.440 ;
        RECT 80.940 161.155 81.110 161.830 ;
        RECT 81.395 161.670 81.565 162.625 ;
        RECT 81.850 162.480 82.020 163.075 ;
        RECT 84.230 162.640 84.690 162.870 ;
        RECT 83.920 162.480 84.090 162.500 ;
        RECT 81.820 161.830 82.050 162.480 ;
        RECT 83.890 161.830 84.120 162.480 ;
        RECT 81.850 161.810 82.020 161.830 ;
        RECT 81.250 161.440 81.710 161.670 ;
        RECT 80.865 160.895 81.185 161.155 ;
        RECT 79.820 159.975 80.140 160.235 ;
        RECT 79.895 159.735 80.065 159.975 ;
        RECT 79.750 159.505 80.210 159.735 ;
        RECT 77.320 158.715 78.140 158.885 ;
        RECT 77.320 158.300 77.550 158.715 ;
        RECT 77.910 158.300 78.140 158.715 ;
        RECT 77.350 158.280 77.520 158.300 ;
        RECT 77.940 158.280 78.110 158.300 ;
        RECT 78.395 158.095 78.565 159.055 ;
        RECT 78.820 158.300 79.050 159.300 ;
        RECT 79.410 158.300 79.640 159.300 ;
        RECT 76.750 157.865 77.210 158.095 ;
        RECT 78.250 157.865 78.710 158.095 ;
        RECT 78.850 157.705 79.020 158.300 ;
        RECT 79.440 158.280 79.610 158.300 ;
        RECT 79.895 158.095 80.065 159.505 ;
        RECT 80.350 159.300 80.520 159.320 ;
        RECT 80.940 159.300 81.110 160.895 ;
        RECT 81.395 159.735 81.565 161.440 ;
        RECT 83.920 160.695 84.090 161.830 ;
        RECT 84.375 161.670 84.545 162.640 ;
        RECT 84.830 162.480 85.000 163.075 ;
        RECT 85.730 162.640 86.190 162.870 ;
        RECT 85.420 162.480 85.590 162.500 ;
        RECT 84.800 161.830 85.030 162.480 ;
        RECT 85.390 161.830 85.620 162.480 ;
        RECT 84.830 161.810 85.000 161.830 ;
        RECT 84.230 161.440 84.690 161.670 ;
        RECT 83.845 160.435 84.165 160.695 ;
        RECT 81.250 159.505 81.710 159.735 ;
        RECT 81.395 159.315 81.565 159.505 ;
        RECT 80.320 158.300 80.550 159.300 ;
        RECT 80.910 158.300 81.140 159.300 ;
        RECT 81.320 159.055 81.640 159.315 ;
        RECT 81.850 159.300 82.020 159.320 ;
        RECT 83.920 159.300 84.090 160.435 ;
        RECT 84.375 160.235 84.545 161.440 ;
        RECT 85.420 160.695 85.590 161.830 ;
        RECT 85.875 161.670 86.045 162.640 ;
        RECT 86.330 162.480 86.500 163.075 ;
        RECT 87.230 162.640 87.690 162.870 ;
        RECT 86.920 162.480 87.090 162.500 ;
        RECT 86.300 161.830 86.530 162.480 ;
        RECT 86.890 161.830 87.120 162.480 ;
        RECT 87.375 162.075 87.545 162.640 ;
        RECT 87.830 162.480 88.000 163.075 ;
        RECT 88.730 162.640 89.190 162.870 ;
        RECT 88.420 162.480 88.590 162.500 ;
        RECT 86.330 161.810 86.500 161.830 ;
        RECT 85.730 161.440 86.190 161.670 ;
        RECT 85.345 160.435 85.665 160.695 ;
        RECT 84.300 159.975 84.620 160.235 ;
        RECT 84.375 159.735 84.545 159.975 ;
        RECT 85.875 159.735 86.045 161.440 ;
        RECT 86.920 160.695 87.090 161.830 ;
        RECT 87.300 161.815 87.620 162.075 ;
        RECT 87.800 161.830 88.030 162.480 ;
        RECT 88.390 161.830 88.620 162.480 ;
        RECT 87.375 161.670 87.545 161.815 ;
        RECT 87.830 161.810 88.000 161.830 ;
        RECT 87.230 161.440 87.690 161.670 ;
        RECT 86.845 160.435 87.165 160.695 ;
        RECT 86.920 160.235 87.090 160.435 ;
        RECT 86.845 159.975 87.165 160.235 ;
        RECT 84.230 159.505 84.690 159.735 ;
        RECT 85.730 159.505 86.190 159.735 ;
        RECT 79.750 157.865 80.210 158.095 ;
        RECT 80.350 157.705 80.520 158.300 ;
        RECT 80.940 158.280 81.110 158.300 ;
        RECT 81.395 158.095 81.565 159.055 ;
        RECT 81.820 158.300 82.050 159.300 ;
        RECT 83.890 158.300 84.120 159.300 ;
        RECT 81.250 157.865 81.710 158.095 ;
        RECT 81.850 157.705 82.020 158.300 ;
        RECT 83.920 158.280 84.090 158.300 ;
        RECT 84.375 158.095 84.545 159.505 ;
        RECT 84.830 159.300 85.000 159.320 ;
        RECT 85.420 159.300 85.590 159.320 ;
        RECT 85.875 159.315 86.045 159.505 ;
        RECT 84.800 158.885 85.030 159.300 ;
        RECT 85.390 158.885 85.620 159.300 ;
        RECT 85.800 159.055 86.120 159.315 ;
        RECT 86.330 159.300 86.500 159.320 ;
        RECT 86.920 159.300 87.090 159.975 ;
        RECT 87.375 159.735 87.545 161.440 ;
        RECT 88.420 160.695 88.590 161.830 ;
        RECT 88.875 161.670 89.045 162.640 ;
        RECT 89.330 162.480 89.500 163.075 ;
        RECT 90.230 162.640 90.690 162.870 ;
        RECT 89.920 162.480 90.090 162.500 ;
        RECT 89.300 161.830 89.530 162.480 ;
        RECT 89.890 161.830 90.120 162.480 ;
        RECT 89.330 161.810 89.500 161.830 ;
        RECT 88.730 161.440 89.190 161.670 ;
        RECT 88.875 161.155 89.045 161.440 ;
        RECT 88.800 160.895 89.120 161.155 ;
        RECT 88.345 160.435 88.665 160.695 ;
        RECT 88.875 159.735 89.045 160.895 ;
        RECT 89.920 160.695 90.090 161.830 ;
        RECT 90.375 161.670 90.545 162.640 ;
        RECT 90.830 162.480 91.000 163.075 ;
        RECT 91.730 162.640 92.190 162.870 ;
        RECT 91.420 162.480 91.590 162.500 ;
        RECT 90.800 161.830 91.030 162.480 ;
        RECT 91.390 161.830 91.620 162.480 ;
        RECT 90.830 161.810 91.000 161.830 ;
        RECT 90.230 161.440 90.690 161.670 ;
        RECT 89.845 160.435 90.165 160.695 ;
        RECT 87.230 159.505 87.690 159.735 ;
        RECT 88.730 159.505 89.190 159.735 ;
        RECT 84.800 158.715 85.620 158.885 ;
        RECT 84.800 158.300 85.030 158.715 ;
        RECT 85.390 158.300 85.620 158.715 ;
        RECT 84.830 158.280 85.000 158.300 ;
        RECT 85.420 158.280 85.590 158.300 ;
        RECT 85.875 158.095 86.045 159.055 ;
        RECT 86.300 158.300 86.530 159.300 ;
        RECT 86.890 158.300 87.120 159.300 ;
        RECT 84.230 157.865 84.690 158.095 ;
        RECT 85.730 157.865 86.190 158.095 ;
        RECT 86.330 157.705 86.500 158.300 ;
        RECT 86.920 158.280 87.090 158.300 ;
        RECT 87.375 158.095 87.545 159.505 ;
        RECT 87.830 159.300 88.000 159.320 ;
        RECT 88.420 159.300 88.590 159.320 ;
        RECT 87.800 158.885 88.030 159.300 ;
        RECT 88.390 158.885 88.620 159.300 ;
        RECT 87.800 158.715 88.620 158.885 ;
        RECT 87.800 158.300 88.030 158.715 ;
        RECT 88.390 158.300 88.620 158.715 ;
        RECT 87.830 158.280 88.000 158.300 ;
        RECT 88.420 158.280 88.590 158.300 ;
        RECT 88.875 158.095 89.045 159.505 ;
        RECT 89.330 159.300 89.500 159.320 ;
        RECT 89.920 159.315 90.090 160.435 ;
        RECT 90.375 160.235 90.545 161.440 ;
        RECT 91.420 160.695 91.590 161.830 ;
        RECT 91.875 161.670 92.045 162.640 ;
        RECT 92.330 162.480 92.500 163.075 ;
        RECT 93.300 162.870 93.620 162.915 ;
        RECT 93.230 162.640 93.690 162.870 ;
        RECT 92.920 162.480 93.090 162.500 ;
        RECT 92.300 161.830 92.530 162.480 ;
        RECT 92.890 162.075 93.120 162.480 ;
        RECT 92.330 161.810 92.500 161.830 ;
        RECT 92.845 161.815 93.165 162.075 ;
        RECT 91.730 161.440 92.190 161.670 ;
        RECT 91.345 160.435 91.665 160.695 ;
        RECT 90.300 159.975 90.620 160.235 ;
        RECT 90.375 159.735 90.545 159.975 ;
        RECT 91.875 159.735 92.045 161.440 ;
        RECT 90.230 159.505 90.690 159.735 ;
        RECT 91.730 159.505 92.190 159.735 ;
        RECT 89.300 158.300 89.530 159.300 ;
        RECT 89.845 159.055 90.165 159.315 ;
        RECT 89.890 158.300 90.120 159.055 ;
        RECT 87.230 157.865 87.690 158.095 ;
        RECT 88.730 157.865 89.190 158.095 ;
        RECT 89.330 157.705 89.500 158.300 ;
        RECT 89.920 158.280 90.090 158.300 ;
        RECT 90.375 158.095 90.545 159.505 ;
        RECT 90.830 159.300 91.000 159.320 ;
        RECT 91.420 159.300 91.590 159.320 ;
        RECT 91.875 159.315 92.045 159.505 ;
        RECT 90.800 158.885 91.030 159.300 ;
        RECT 91.390 158.885 91.620 159.300 ;
        RECT 91.800 159.055 92.120 159.315 ;
        RECT 92.330 159.300 92.500 159.320 ;
        RECT 92.920 159.300 93.090 161.815 ;
        RECT 93.375 161.670 93.545 162.640 ;
        RECT 93.830 162.480 94.000 163.075 ;
        RECT 94.800 162.870 95.120 162.885 ;
        RECT 94.730 162.640 95.190 162.870 ;
        RECT 94.800 162.625 95.120 162.640 ;
        RECT 94.420 162.480 94.590 162.500 ;
        RECT 93.800 161.830 94.030 162.480 ;
        RECT 94.390 161.830 94.620 162.480 ;
        RECT 93.830 161.810 94.000 161.830 ;
        RECT 93.230 161.440 93.690 161.670 ;
        RECT 93.375 160.235 93.545 161.440 ;
        RECT 94.420 161.155 94.590 161.830 ;
        RECT 94.875 161.670 95.045 162.625 ;
        RECT 95.330 162.480 95.500 163.075 ;
        RECT 103.685 163.040 103.985 163.075 ;
        RECT 95.300 161.830 95.530 162.480 ;
        RECT 95.330 161.810 95.500 161.830 ;
        RECT 94.730 161.440 95.190 161.670 ;
        RECT 94.345 160.895 94.665 161.155 ;
        RECT 93.300 159.975 93.620 160.235 ;
        RECT 93.375 159.735 93.545 159.975 ;
        RECT 93.230 159.505 93.690 159.735 ;
        RECT 90.800 158.715 91.620 158.885 ;
        RECT 90.800 158.300 91.030 158.715 ;
        RECT 91.390 158.300 91.620 158.715 ;
        RECT 90.830 158.280 91.000 158.300 ;
        RECT 91.420 158.280 91.590 158.300 ;
        RECT 91.875 158.095 92.045 159.055 ;
        RECT 92.300 158.300 92.530 159.300 ;
        RECT 92.890 158.300 93.120 159.300 ;
        RECT 90.230 157.865 90.690 158.095 ;
        RECT 91.730 157.865 92.190 158.095 ;
        RECT 92.330 157.705 92.500 158.300 ;
        RECT 92.920 158.280 93.090 158.300 ;
        RECT 93.375 158.095 93.545 159.505 ;
        RECT 93.830 159.300 94.000 159.320 ;
        RECT 94.420 159.300 94.590 160.895 ;
        RECT 94.875 159.735 95.045 161.440 ;
        RECT 94.730 159.505 95.190 159.735 ;
        RECT 94.875 159.315 95.045 159.505 ;
        RECT 93.800 158.300 94.030 159.300 ;
        RECT 94.390 158.300 94.620 159.300 ;
        RECT 94.800 159.055 95.120 159.315 ;
        RECT 95.330 159.300 95.500 159.320 ;
        RECT 93.230 157.865 93.690 158.095 ;
        RECT 93.830 157.705 94.000 158.300 ;
        RECT 94.420 158.280 94.590 158.300 ;
        RECT 94.875 158.095 95.045 159.055 ;
        RECT 95.300 158.300 95.530 159.300 ;
        RECT 94.730 157.865 95.190 158.095 ;
        RECT 95.330 157.705 95.500 158.300 ;
        RECT 105.185 157.705 105.485 157.740 ;
        RECT 33.145 157.415 105.485 157.705 ;
        RECT 33.145 157.380 33.445 157.415 ;
        RECT 105.185 157.380 105.485 157.415 ;
        RECT 49.890 156.930 50.150 157.020 ;
        RECT 58.175 156.930 58.435 157.020 ;
        RECT 76.850 156.930 77.110 157.050 ;
        RECT 90.330 156.930 90.590 157.005 ;
        RECT 49.890 156.760 90.590 156.930 ;
        RECT 49.890 156.700 50.150 156.760 ;
        RECT 58.175 156.700 58.435 156.760 ;
        RECT 76.850 156.730 77.110 156.760 ;
        RECT 90.330 156.685 90.590 156.760 ;
        RECT 52.235 156.205 52.495 156.280 ;
        RECT 65.655 156.205 65.915 156.280 ;
        RECT 79.075 156.205 79.335 156.280 ;
        RECT 92.495 156.205 92.755 156.280 ;
        RECT 52.235 156.035 92.755 156.205 ;
        RECT 52.235 155.960 52.495 156.035 ;
        RECT 65.655 155.960 65.915 156.035 ;
        RECT 79.075 155.960 79.335 156.035 ;
        RECT 92.495 155.960 92.755 156.035 ;
        RECT 42.300 155.820 42.560 155.895 ;
        RECT 50.430 155.820 50.690 155.895 ;
        RECT 42.300 155.650 50.690 155.820 ;
        RECT 42.300 155.575 42.560 155.650 ;
        RECT 50.430 155.575 50.690 155.650 ;
        RECT 58.945 155.820 59.205 155.895 ;
        RECT 72.335 155.820 72.655 155.865 ;
        RECT 85.785 155.820 86.045 155.895 ;
        RECT 99.205 155.820 99.465 155.895 ;
        RECT 58.945 155.650 99.465 155.820 ;
        RECT 58.945 155.575 59.205 155.650 ;
        RECT 72.335 155.605 72.655 155.650 ;
        RECT 85.785 155.575 86.045 155.650 ;
        RECT 99.205 155.575 99.465 155.650 ;
        RECT 39.235 155.435 39.495 155.510 ;
        RECT 63.850 155.435 64.110 155.510 ;
        RECT 39.235 155.265 64.110 155.435 ;
        RECT 39.235 155.190 39.495 155.265 ;
        RECT 63.850 155.190 64.110 155.265 ;
        RECT 49.010 155.050 49.270 155.125 ;
        RECT 77.270 155.050 77.530 155.125 ;
        RECT 49.010 154.880 77.530 155.050 ;
        RECT 49.010 154.805 49.270 154.880 ;
        RECT 77.270 154.805 77.530 154.880 ;
        RECT 45.945 154.665 46.205 154.740 ;
        RECT 90.690 154.665 90.950 154.740 ;
        RECT 45.945 154.495 90.950 154.665 ;
        RECT 45.945 154.420 46.205 154.495 ;
        RECT 90.690 154.420 90.950 154.495 ;
        RECT 36.145 154.115 36.435 154.325 ;
        RECT 37.030 154.115 37.680 154.145 ;
        RECT 40.210 154.115 41.210 154.145 ;
        RECT 41.805 154.115 42.095 154.325 ;
        RECT 36.145 153.945 37.700 154.115 ;
        RECT 40.190 154.050 42.095 154.115 ;
        RECT 42.855 154.115 43.145 154.325 ;
        RECT 43.740 154.115 44.390 154.145 ;
        RECT 46.920 154.115 47.920 154.145 ;
        RECT 48.515 154.115 48.805 154.325 ;
        RECT 40.190 153.945 42.100 154.050 ;
        RECT 36.145 152.615 36.435 153.945 ;
        RECT 37.030 153.915 37.680 153.945 ;
        RECT 40.210 153.915 41.210 153.945 ;
        RECT 36.640 153.660 36.870 153.805 ;
        RECT 37.010 153.660 37.270 153.735 ;
        RECT 37.840 153.660 38.070 153.805 ;
        RECT 39.775 153.660 40.005 153.805 ;
        RECT 41.415 153.660 41.645 153.805 ;
        RECT 41.800 153.690 42.100 153.945 ;
        RECT 42.855 153.945 44.410 154.115 ;
        RECT 46.900 154.050 48.805 154.115 ;
        RECT 49.565 154.115 49.855 154.325 ;
        RECT 50.450 154.115 51.100 154.145 ;
        RECT 53.630 154.115 54.630 154.145 ;
        RECT 55.225 154.115 55.515 154.325 ;
        RECT 46.900 153.945 48.810 154.050 ;
        RECT 36.640 153.490 41.645 153.660 ;
        RECT 36.640 153.345 36.870 153.490 ;
        RECT 37.010 153.415 37.270 153.490 ;
        RECT 37.840 153.345 38.070 153.490 ;
        RECT 39.775 153.345 40.005 153.490 ;
        RECT 41.415 153.345 41.645 153.490 ;
        RECT 40.970 153.235 41.230 153.280 ;
        RECT 37.030 153.205 37.680 153.235 ;
        RECT 40.210 153.205 41.230 153.235 ;
        RECT 37.010 153.035 41.230 153.205 ;
        RECT 37.030 153.005 37.680 153.035 ;
        RECT 40.210 153.005 41.230 153.035 ;
        RECT 40.970 152.960 41.230 153.005 ;
        RECT 37.030 152.615 37.680 152.645 ;
        RECT 40.210 152.615 41.210 152.645 ;
        RECT 41.805 152.615 42.095 153.690 ;
        RECT 36.145 152.550 37.700 152.615 ;
        RECT 36.140 152.445 37.700 152.550 ;
        RECT 40.190 152.445 42.095 152.615 ;
        RECT 42.855 153.660 43.145 153.945 ;
        RECT 43.740 153.915 44.390 153.945 ;
        RECT 46.920 153.915 47.920 153.945 ;
        RECT 43.350 153.660 43.580 153.805 ;
        RECT 44.550 153.660 44.780 153.805 ;
        RECT 46.485 153.660 46.715 153.805 ;
        RECT 48.125 153.660 48.355 153.805 ;
        RECT 48.510 153.690 48.810 153.945 ;
        RECT 49.565 153.945 51.120 154.115 ;
        RECT 53.610 154.050 55.515 154.115 ;
        RECT 56.275 154.115 56.565 154.325 ;
        RECT 57.160 154.115 57.810 154.145 ;
        RECT 60.340 154.115 61.340 154.145 ;
        RECT 61.935 154.115 62.225 154.325 ;
        RECT 53.610 153.945 55.520 154.050 ;
        RECT 42.855 153.490 48.355 153.660 ;
        RECT 42.855 152.615 43.145 153.490 ;
        RECT 43.350 153.345 43.580 153.490 ;
        RECT 44.550 153.345 44.780 153.490 ;
        RECT 46.485 153.345 46.715 153.490 ;
        RECT 48.125 153.345 48.355 153.490 ;
        RECT 43.740 153.205 44.390 153.235 ;
        RECT 46.920 153.205 47.920 153.235 ;
        RECT 43.720 153.035 47.940 153.205 ;
        RECT 43.740 153.005 44.390 153.035 ;
        RECT 46.920 153.005 47.920 153.035 ;
        RECT 43.740 152.615 44.390 152.645 ;
        RECT 46.920 152.615 47.920 152.645 ;
        RECT 48.515 152.615 48.805 153.690 ;
        RECT 42.855 152.550 44.410 152.615 ;
        RECT 36.140 152.190 36.440 152.445 ;
        RECT 37.030 152.415 37.680 152.445 ;
        RECT 40.210 152.415 41.210 152.445 ;
        RECT 36.145 151.115 36.435 152.190 ;
        RECT 36.640 152.160 36.870 152.305 ;
        RECT 37.840 152.160 38.070 152.305 ;
        RECT 38.785 152.160 39.105 152.205 ;
        RECT 39.775 152.160 40.005 152.305 ;
        RECT 41.415 152.160 41.645 152.305 ;
        RECT 36.640 151.990 41.645 152.160 ;
        RECT 36.640 151.845 36.870 151.990 ;
        RECT 37.840 151.845 38.070 151.990 ;
        RECT 38.785 151.945 39.105 151.990 ;
        RECT 39.775 151.845 40.005 151.990 ;
        RECT 41.415 151.845 41.645 151.990 ;
        RECT 37.030 151.705 37.680 151.735 ;
        RECT 38.815 151.705 39.075 151.780 ;
        RECT 40.130 151.735 40.390 151.780 ;
        RECT 40.130 151.705 41.210 151.735 ;
        RECT 37.010 151.535 41.230 151.705 ;
        RECT 37.030 151.505 37.680 151.535 ;
        RECT 38.815 151.460 39.075 151.535 ;
        RECT 40.130 151.505 41.210 151.535 ;
        RECT 40.130 151.460 40.390 151.505 ;
        RECT 37.030 151.115 37.680 151.145 ;
        RECT 40.210 151.115 41.210 151.145 ;
        RECT 41.805 151.115 42.095 152.445 ;
        RECT 42.850 152.445 44.410 152.550 ;
        RECT 46.900 152.445 48.805 152.615 ;
        RECT 49.565 152.615 49.855 153.945 ;
        RECT 50.450 153.915 51.100 153.945 ;
        RECT 53.630 153.915 54.630 153.945 ;
        RECT 50.060 153.660 50.290 153.805 ;
        RECT 50.430 153.660 50.690 153.735 ;
        RECT 51.260 153.660 51.490 153.805 ;
        RECT 53.195 153.660 53.425 153.805 ;
        RECT 54.835 153.660 55.065 153.805 ;
        RECT 55.220 153.690 55.520 153.945 ;
        RECT 56.275 153.945 57.830 154.115 ;
        RECT 60.320 154.050 62.225 154.115 ;
        RECT 62.985 154.115 63.275 154.325 ;
        RECT 63.870 154.115 64.520 154.145 ;
        RECT 67.050 154.115 68.050 154.145 ;
        RECT 68.645 154.115 68.935 154.325 ;
        RECT 60.320 153.945 62.230 154.050 ;
        RECT 50.060 153.490 55.065 153.660 ;
        RECT 50.060 153.345 50.290 153.490 ;
        RECT 50.430 153.415 50.690 153.490 ;
        RECT 51.260 153.345 51.490 153.490 ;
        RECT 53.195 153.345 53.425 153.490 ;
        RECT 54.835 153.345 55.065 153.490 ;
        RECT 54.390 153.235 54.650 153.280 ;
        RECT 50.450 153.205 51.100 153.235 ;
        RECT 53.630 153.205 54.650 153.235 ;
        RECT 50.430 153.035 54.650 153.205 ;
        RECT 50.450 153.005 51.100 153.035 ;
        RECT 53.630 153.005 54.650 153.035 ;
        RECT 54.390 152.960 54.650 153.005 ;
        RECT 50.450 152.615 51.100 152.645 ;
        RECT 53.630 152.615 54.630 152.645 ;
        RECT 55.225 152.615 55.515 153.690 ;
        RECT 49.565 152.550 51.120 152.615 ;
        RECT 42.850 152.190 43.150 152.445 ;
        RECT 43.740 152.415 44.390 152.445 ;
        RECT 46.920 152.415 47.920 152.445 ;
        RECT 36.145 150.945 37.700 151.115 ;
        RECT 40.190 151.050 42.095 151.115 ;
        RECT 42.855 151.115 43.145 152.190 ;
        RECT 43.350 152.160 43.580 152.305 ;
        RECT 44.550 152.160 44.780 152.305 ;
        RECT 45.495 152.160 45.815 152.205 ;
        RECT 46.485 152.160 46.715 152.305 ;
        RECT 48.125 152.160 48.355 152.305 ;
        RECT 43.350 151.990 48.355 152.160 ;
        RECT 43.350 151.845 43.580 151.990 ;
        RECT 44.550 151.845 44.780 151.990 ;
        RECT 45.495 151.945 45.815 151.990 ;
        RECT 46.485 151.845 46.715 151.990 ;
        RECT 48.125 151.845 48.355 151.990 ;
        RECT 43.740 151.705 44.390 151.735 ;
        RECT 45.525 151.705 45.785 151.780 ;
        RECT 46.920 151.705 47.920 151.735 ;
        RECT 43.720 151.535 47.940 151.705 ;
        RECT 43.740 151.505 44.390 151.535 ;
        RECT 45.525 151.460 45.785 151.535 ;
        RECT 46.460 151.375 46.630 151.535 ;
        RECT 46.920 151.505 47.920 151.535 ;
        RECT 43.740 151.115 44.390 151.145 ;
        RECT 40.190 150.945 42.100 151.050 ;
        RECT 36.145 149.615 36.435 150.945 ;
        RECT 37.030 150.915 37.680 150.945 ;
        RECT 40.210 150.915 41.210 150.945 ;
        RECT 36.640 150.660 36.870 150.805 ;
        RECT 37.840 150.660 38.070 150.805 ;
        RECT 38.815 150.660 39.075 150.735 ;
        RECT 39.775 150.660 40.005 150.805 ;
        RECT 41.415 150.660 41.645 150.805 ;
        RECT 41.800 150.690 42.100 150.945 ;
        RECT 42.855 150.945 44.410 151.115 ;
        RECT 46.415 151.055 46.675 151.375 ;
        RECT 46.920 151.115 47.920 151.145 ;
        RECT 48.515 151.115 48.805 152.445 ;
        RECT 49.560 152.445 51.120 152.550 ;
        RECT 53.610 152.445 55.515 152.615 ;
        RECT 56.275 153.660 56.565 153.945 ;
        RECT 57.160 153.915 57.810 153.945 ;
        RECT 60.340 153.915 61.340 153.945 ;
        RECT 56.770 153.660 57.000 153.805 ;
        RECT 57.970 153.660 58.200 153.805 ;
        RECT 59.905 153.660 60.135 153.805 ;
        RECT 61.545 153.660 61.775 153.805 ;
        RECT 61.930 153.690 62.230 153.945 ;
        RECT 62.985 153.945 64.540 154.115 ;
        RECT 67.030 154.050 68.935 154.115 ;
        RECT 69.695 154.115 69.985 154.325 ;
        RECT 70.580 154.115 71.230 154.145 ;
        RECT 73.760 154.115 74.760 154.145 ;
        RECT 75.355 154.115 75.645 154.325 ;
        RECT 67.030 153.945 68.940 154.050 ;
        RECT 56.275 153.490 61.775 153.660 ;
        RECT 56.275 152.615 56.565 153.490 ;
        RECT 56.770 153.345 57.000 153.490 ;
        RECT 57.970 153.345 58.200 153.490 ;
        RECT 59.905 153.345 60.135 153.490 ;
        RECT 61.545 153.345 61.775 153.490 ;
        RECT 57.160 153.205 57.810 153.235 ;
        RECT 60.340 153.205 61.340 153.235 ;
        RECT 57.140 153.035 61.360 153.205 ;
        RECT 57.160 153.005 57.810 153.035 ;
        RECT 60.340 153.005 61.340 153.035 ;
        RECT 57.160 152.615 57.810 152.645 ;
        RECT 60.340 152.615 61.340 152.645 ;
        RECT 61.935 152.615 62.225 153.690 ;
        RECT 56.275 152.550 57.830 152.615 ;
        RECT 49.560 152.190 49.860 152.445 ;
        RECT 50.450 152.415 51.100 152.445 ;
        RECT 53.630 152.415 54.630 152.445 ;
        RECT 46.900 151.050 48.805 151.115 ;
        RECT 49.565 151.115 49.855 152.190 ;
        RECT 50.060 152.160 50.290 152.305 ;
        RECT 51.260 152.160 51.490 152.305 ;
        RECT 52.205 152.160 52.525 152.205 ;
        RECT 53.195 152.160 53.425 152.305 ;
        RECT 54.835 152.160 55.065 152.305 ;
        RECT 50.060 151.990 55.065 152.160 ;
        RECT 50.060 151.845 50.290 151.990 ;
        RECT 51.260 151.845 51.490 151.990 ;
        RECT 52.205 151.945 52.525 151.990 ;
        RECT 53.195 151.845 53.425 151.990 ;
        RECT 54.835 151.845 55.065 151.990 ;
        RECT 50.450 151.705 51.100 151.735 ;
        RECT 52.235 151.705 52.495 151.780 ;
        RECT 53.550 151.735 53.810 151.780 ;
        RECT 53.550 151.705 54.630 151.735 ;
        RECT 50.430 151.535 54.650 151.705 ;
        RECT 50.450 151.505 51.100 151.535 ;
        RECT 52.235 151.460 52.495 151.535 ;
        RECT 53.550 151.505 54.630 151.535 ;
        RECT 53.550 151.460 53.810 151.505 ;
        RECT 50.450 151.115 51.100 151.145 ;
        RECT 53.630 151.115 54.630 151.145 ;
        RECT 55.225 151.115 55.515 152.445 ;
        RECT 56.270 152.445 57.830 152.550 ;
        RECT 60.320 152.445 62.225 152.615 ;
        RECT 62.985 152.615 63.275 153.945 ;
        RECT 63.870 153.915 64.520 153.945 ;
        RECT 67.050 153.915 68.050 153.945 ;
        RECT 63.480 153.660 63.710 153.805 ;
        RECT 63.850 153.660 64.110 153.735 ;
        RECT 64.680 153.660 64.910 153.805 ;
        RECT 66.615 153.660 66.845 153.805 ;
        RECT 68.255 153.660 68.485 153.805 ;
        RECT 68.640 153.690 68.940 153.945 ;
        RECT 69.695 153.945 71.250 154.115 ;
        RECT 73.740 154.050 75.645 154.115 ;
        RECT 76.405 154.115 76.695 154.325 ;
        RECT 77.290 154.115 77.940 154.145 ;
        RECT 80.470 154.115 81.470 154.145 ;
        RECT 82.065 154.115 82.355 154.325 ;
        RECT 73.740 153.945 75.650 154.050 ;
        RECT 63.480 153.490 68.485 153.660 ;
        RECT 63.480 153.345 63.710 153.490 ;
        RECT 63.850 153.415 64.110 153.490 ;
        RECT 64.680 153.345 64.910 153.490 ;
        RECT 66.615 153.345 66.845 153.490 ;
        RECT 68.255 153.345 68.485 153.490 ;
        RECT 67.810 153.235 68.070 153.280 ;
        RECT 63.870 153.205 64.520 153.235 ;
        RECT 67.050 153.205 68.070 153.235 ;
        RECT 63.850 153.035 68.070 153.205 ;
        RECT 63.870 153.005 64.520 153.035 ;
        RECT 67.050 153.005 68.070 153.035 ;
        RECT 67.810 152.960 68.070 153.005 ;
        RECT 63.870 152.615 64.520 152.645 ;
        RECT 67.050 152.615 68.050 152.645 ;
        RECT 68.645 152.615 68.935 153.690 ;
        RECT 62.985 152.550 64.540 152.615 ;
        RECT 56.270 152.190 56.570 152.445 ;
        RECT 57.160 152.415 57.810 152.445 ;
        RECT 60.340 152.415 61.340 152.445 ;
        RECT 46.900 150.945 48.810 151.050 ;
        RECT 36.640 150.490 41.645 150.660 ;
        RECT 36.640 150.345 36.870 150.490 ;
        RECT 37.840 150.345 38.070 150.490 ;
        RECT 38.815 150.415 39.075 150.490 ;
        RECT 39.775 150.345 40.005 150.490 ;
        RECT 41.415 150.345 41.645 150.490 ;
        RECT 40.550 150.235 40.810 150.280 ;
        RECT 37.030 150.205 37.680 150.235 ;
        RECT 40.210 150.205 41.210 150.235 ;
        RECT 37.010 150.035 41.230 150.205 ;
        RECT 37.030 150.005 37.680 150.035 ;
        RECT 40.210 150.005 41.210 150.035 ;
        RECT 40.550 149.960 40.810 150.005 ;
        RECT 37.030 149.615 37.680 149.645 ;
        RECT 40.210 149.615 41.210 149.645 ;
        RECT 41.805 149.615 42.095 150.690 ;
        RECT 36.145 149.550 37.700 149.615 ;
        RECT 36.140 149.445 37.700 149.550 ;
        RECT 40.190 149.445 42.095 149.615 ;
        RECT 42.855 149.615 43.145 150.945 ;
        RECT 43.740 150.915 44.390 150.945 ;
        RECT 46.920 150.915 47.920 150.945 ;
        RECT 43.350 150.660 43.580 150.805 ;
        RECT 44.550 150.660 44.780 150.805 ;
        RECT 45.525 150.660 45.785 150.735 ;
        RECT 46.485 150.660 46.715 150.805 ;
        RECT 48.125 150.660 48.355 150.805 ;
        RECT 48.510 150.690 48.810 150.945 ;
        RECT 49.565 150.945 51.120 151.115 ;
        RECT 53.610 151.050 55.515 151.115 ;
        RECT 56.275 151.115 56.565 152.190 ;
        RECT 56.770 152.160 57.000 152.305 ;
        RECT 57.970 152.160 58.200 152.305 ;
        RECT 58.915 152.160 59.235 152.205 ;
        RECT 59.905 152.160 60.135 152.305 ;
        RECT 61.545 152.160 61.775 152.305 ;
        RECT 56.770 151.990 61.775 152.160 ;
        RECT 56.770 151.845 57.000 151.990 ;
        RECT 57.970 151.845 58.200 151.990 ;
        RECT 58.915 151.945 59.235 151.990 ;
        RECT 59.905 151.845 60.135 151.990 ;
        RECT 61.545 151.845 61.775 151.990 ;
        RECT 57.160 151.705 57.810 151.735 ;
        RECT 58.945 151.705 59.205 151.780 ;
        RECT 60.340 151.705 61.340 151.735 ;
        RECT 57.140 151.535 61.360 151.705 ;
        RECT 57.160 151.505 57.810 151.535 ;
        RECT 58.945 151.460 59.205 151.535 ;
        RECT 59.880 151.375 60.050 151.535 ;
        RECT 60.340 151.505 61.340 151.535 ;
        RECT 57.160 151.115 57.810 151.145 ;
        RECT 53.610 150.945 55.520 151.050 ;
        RECT 43.350 150.490 48.355 150.660 ;
        RECT 43.350 150.345 43.580 150.490 ;
        RECT 44.550 150.345 44.780 150.490 ;
        RECT 45.525 150.415 45.785 150.490 ;
        RECT 46.485 150.345 46.715 150.490 ;
        RECT 48.125 150.345 48.355 150.490 ;
        RECT 43.720 150.235 43.980 150.280 ;
        RECT 43.720 150.205 44.390 150.235 ;
        RECT 46.920 150.205 47.920 150.235 ;
        RECT 43.720 150.035 47.940 150.205 ;
        RECT 43.720 150.005 44.390 150.035 ;
        RECT 46.920 150.005 47.920 150.035 ;
        RECT 43.720 149.960 43.980 150.005 ;
        RECT 43.740 149.615 44.390 149.645 ;
        RECT 46.920 149.615 47.920 149.645 ;
        RECT 48.515 149.615 48.805 150.690 ;
        RECT 42.855 149.550 44.410 149.615 ;
        RECT 36.140 149.190 36.440 149.445 ;
        RECT 37.030 149.415 37.680 149.445 ;
        RECT 40.210 149.415 41.210 149.445 ;
        RECT 36.145 148.115 36.435 149.190 ;
        RECT 36.640 149.160 36.870 149.305 ;
        RECT 37.840 149.160 38.070 149.305 ;
        RECT 39.775 149.235 40.005 149.305 ;
        RECT 39.710 149.160 40.005 149.235 ;
        RECT 41.415 149.160 41.645 149.305 ;
        RECT 36.640 148.990 41.645 149.160 ;
        RECT 36.640 148.845 36.870 148.990 ;
        RECT 37.840 148.845 38.070 148.990 ;
        RECT 39.710 148.915 40.005 148.990 ;
        RECT 39.775 148.845 40.005 148.915 ;
        RECT 41.415 148.845 41.645 148.990 ;
        RECT 37.030 148.705 37.680 148.735 ;
        RECT 38.815 148.705 39.075 148.780 ;
        RECT 40.210 148.705 41.210 148.735 ;
        RECT 37.010 148.535 39.075 148.705 ;
        RECT 40.190 148.535 41.230 148.705 ;
        RECT 37.030 148.505 37.680 148.535 ;
        RECT 38.815 148.460 39.075 148.535 ;
        RECT 40.210 148.505 41.210 148.535 ;
        RECT 40.625 148.145 40.795 148.505 ;
        RECT 37.030 148.115 37.680 148.145 ;
        RECT 40.210 148.115 41.210 148.145 ;
        RECT 36.145 147.945 37.700 148.115 ;
        RECT 40.190 147.945 41.230 148.115 ;
        RECT 41.805 148.050 42.095 149.445 ;
        RECT 42.850 149.445 44.410 149.550 ;
        RECT 46.900 149.445 48.805 149.615 ;
        RECT 49.565 149.615 49.855 150.945 ;
        RECT 50.450 150.915 51.100 150.945 ;
        RECT 53.630 150.915 54.630 150.945 ;
        RECT 50.060 150.660 50.290 150.805 ;
        RECT 51.260 150.660 51.490 150.805 ;
        RECT 52.235 150.660 52.495 150.735 ;
        RECT 53.195 150.660 53.425 150.805 ;
        RECT 54.835 150.660 55.065 150.805 ;
        RECT 55.220 150.690 55.520 150.945 ;
        RECT 56.275 150.945 57.830 151.115 ;
        RECT 59.835 151.055 60.095 151.375 ;
        RECT 60.340 151.115 61.340 151.145 ;
        RECT 61.935 151.115 62.225 152.445 ;
        RECT 62.980 152.445 64.540 152.550 ;
        RECT 67.030 152.445 68.935 152.615 ;
        RECT 69.695 153.660 69.985 153.945 ;
        RECT 70.580 153.915 71.230 153.945 ;
        RECT 73.760 153.915 74.760 153.945 ;
        RECT 70.190 153.660 70.420 153.805 ;
        RECT 71.390 153.660 71.620 153.805 ;
        RECT 73.325 153.660 73.555 153.805 ;
        RECT 74.965 153.660 75.195 153.805 ;
        RECT 75.350 153.690 75.650 153.945 ;
        RECT 76.405 153.945 77.960 154.115 ;
        RECT 80.450 154.050 82.355 154.115 ;
        RECT 83.115 154.115 83.405 154.325 ;
        RECT 84.000 154.115 84.650 154.145 ;
        RECT 87.180 154.115 88.180 154.145 ;
        RECT 88.775 154.115 89.065 154.325 ;
        RECT 80.450 153.945 82.360 154.050 ;
        RECT 69.695 153.490 75.195 153.660 ;
        RECT 69.695 152.615 69.985 153.490 ;
        RECT 70.190 153.345 70.420 153.490 ;
        RECT 71.390 153.345 71.620 153.490 ;
        RECT 73.325 153.345 73.555 153.490 ;
        RECT 74.965 153.345 75.195 153.490 ;
        RECT 70.580 153.205 71.230 153.235 ;
        RECT 73.760 153.205 74.760 153.235 ;
        RECT 70.560 153.035 74.780 153.205 ;
        RECT 70.580 153.005 71.230 153.035 ;
        RECT 73.760 153.005 74.760 153.035 ;
        RECT 70.580 152.615 71.230 152.645 ;
        RECT 73.760 152.615 74.760 152.645 ;
        RECT 75.355 152.615 75.645 153.690 ;
        RECT 69.695 152.550 71.250 152.615 ;
        RECT 62.980 152.190 63.280 152.445 ;
        RECT 63.870 152.415 64.520 152.445 ;
        RECT 67.050 152.415 68.050 152.445 ;
        RECT 60.320 151.050 62.225 151.115 ;
        RECT 62.985 151.115 63.275 152.190 ;
        RECT 63.480 152.160 63.710 152.305 ;
        RECT 64.680 152.160 64.910 152.305 ;
        RECT 65.625 152.160 65.945 152.205 ;
        RECT 66.615 152.160 66.845 152.305 ;
        RECT 68.255 152.160 68.485 152.305 ;
        RECT 63.480 151.990 68.485 152.160 ;
        RECT 63.480 151.845 63.710 151.990 ;
        RECT 64.680 151.845 64.910 151.990 ;
        RECT 65.625 151.945 65.945 151.990 ;
        RECT 66.615 151.845 66.845 151.990 ;
        RECT 68.255 151.845 68.485 151.990 ;
        RECT 63.870 151.705 64.520 151.735 ;
        RECT 65.655 151.705 65.915 151.780 ;
        RECT 66.970 151.735 67.230 151.780 ;
        RECT 66.970 151.705 68.050 151.735 ;
        RECT 63.850 151.535 68.070 151.705 ;
        RECT 63.870 151.505 64.520 151.535 ;
        RECT 65.655 151.460 65.915 151.535 ;
        RECT 66.970 151.505 68.050 151.535 ;
        RECT 66.970 151.460 67.230 151.505 ;
        RECT 63.870 151.115 64.520 151.145 ;
        RECT 67.050 151.115 68.050 151.145 ;
        RECT 68.645 151.115 68.935 152.445 ;
        RECT 69.690 152.445 71.250 152.550 ;
        RECT 73.740 152.445 75.645 152.615 ;
        RECT 76.405 152.615 76.695 153.945 ;
        RECT 77.290 153.915 77.940 153.945 ;
        RECT 80.470 153.915 81.470 153.945 ;
        RECT 76.900 153.660 77.130 153.805 ;
        RECT 77.270 153.660 77.530 153.735 ;
        RECT 78.100 153.660 78.330 153.805 ;
        RECT 80.035 153.660 80.265 153.805 ;
        RECT 81.675 153.660 81.905 153.805 ;
        RECT 82.060 153.690 82.360 153.945 ;
        RECT 83.115 153.945 84.670 154.115 ;
        RECT 87.160 154.050 89.065 154.115 ;
        RECT 89.825 154.115 90.115 154.325 ;
        RECT 90.710 154.115 91.360 154.145 ;
        RECT 93.890 154.115 94.890 154.145 ;
        RECT 95.485 154.115 95.775 154.325 ;
        RECT 87.160 153.945 89.070 154.050 ;
        RECT 76.900 153.490 81.905 153.660 ;
        RECT 76.900 153.345 77.130 153.490 ;
        RECT 77.270 153.415 77.530 153.490 ;
        RECT 78.100 153.345 78.330 153.490 ;
        RECT 80.035 153.345 80.265 153.490 ;
        RECT 81.675 153.345 81.905 153.490 ;
        RECT 81.230 153.235 81.490 153.280 ;
        RECT 77.290 153.205 77.940 153.235 ;
        RECT 80.470 153.205 81.490 153.235 ;
        RECT 77.270 153.035 81.490 153.205 ;
        RECT 77.290 153.005 77.940 153.035 ;
        RECT 80.470 153.005 81.490 153.035 ;
        RECT 81.230 152.960 81.490 153.005 ;
        RECT 77.290 152.615 77.940 152.645 ;
        RECT 80.470 152.615 81.470 152.645 ;
        RECT 82.065 152.615 82.355 153.690 ;
        RECT 76.405 152.550 77.960 152.615 ;
        RECT 69.690 152.190 69.990 152.445 ;
        RECT 70.580 152.415 71.230 152.445 ;
        RECT 73.760 152.415 74.760 152.445 ;
        RECT 60.320 150.945 62.230 151.050 ;
        RECT 50.060 150.490 55.065 150.660 ;
        RECT 50.060 150.345 50.290 150.490 ;
        RECT 51.260 150.345 51.490 150.490 ;
        RECT 52.235 150.415 52.495 150.490 ;
        RECT 53.195 150.345 53.425 150.490 ;
        RECT 54.835 150.345 55.065 150.490 ;
        RECT 53.970 150.235 54.230 150.280 ;
        RECT 50.450 150.205 51.100 150.235 ;
        RECT 53.630 150.205 54.630 150.235 ;
        RECT 50.430 150.035 54.650 150.205 ;
        RECT 50.450 150.005 51.100 150.035 ;
        RECT 53.630 150.005 54.630 150.035 ;
        RECT 53.970 149.960 54.230 150.005 ;
        RECT 50.450 149.615 51.100 149.645 ;
        RECT 53.630 149.615 54.630 149.645 ;
        RECT 55.225 149.615 55.515 150.690 ;
        RECT 49.565 149.550 51.120 149.615 ;
        RECT 42.850 149.190 43.150 149.445 ;
        RECT 43.740 149.415 44.390 149.445 ;
        RECT 46.920 149.415 47.920 149.445 ;
        RECT 42.855 148.115 43.145 149.190 ;
        RECT 43.350 149.160 43.580 149.305 ;
        RECT 44.550 149.160 44.780 149.305 ;
        RECT 46.485 149.235 46.715 149.305 ;
        RECT 46.420 149.160 46.715 149.235 ;
        RECT 48.125 149.160 48.355 149.305 ;
        RECT 43.350 148.990 48.355 149.160 ;
        RECT 43.350 148.845 43.580 148.990 ;
        RECT 44.550 148.845 44.780 148.990 ;
        RECT 46.420 148.915 46.715 148.990 ;
        RECT 46.485 148.845 46.715 148.915 ;
        RECT 48.125 148.845 48.355 148.990 ;
        RECT 43.740 148.705 44.390 148.735 ;
        RECT 45.525 148.705 45.785 148.780 ;
        RECT 46.920 148.705 47.920 148.735 ;
        RECT 43.720 148.535 45.785 148.705 ;
        RECT 46.900 148.535 47.940 148.705 ;
        RECT 43.740 148.505 44.390 148.535 ;
        RECT 45.525 148.460 45.785 148.535 ;
        RECT 46.920 148.505 47.920 148.535 ;
        RECT 47.335 148.145 47.505 148.505 ;
        RECT 43.740 148.115 44.390 148.145 ;
        RECT 46.920 148.115 47.920 148.145 ;
        RECT 36.145 146.615 36.435 147.945 ;
        RECT 37.030 147.915 37.680 147.945 ;
        RECT 40.210 147.915 41.210 147.945 ;
        RECT 36.640 147.660 36.870 147.805 ;
        RECT 37.840 147.660 38.070 147.805 ;
        RECT 39.775 147.660 40.005 147.805 ;
        RECT 40.550 147.660 40.810 147.735 ;
        RECT 41.415 147.660 41.645 147.805 ;
        RECT 41.800 147.690 42.100 148.050 ;
        RECT 42.855 147.945 44.410 148.115 ;
        RECT 46.900 147.945 47.940 148.115 ;
        RECT 48.515 148.050 48.805 149.445 ;
        RECT 49.560 149.445 51.120 149.550 ;
        RECT 53.610 149.445 55.515 149.615 ;
        RECT 56.275 149.615 56.565 150.945 ;
        RECT 57.160 150.915 57.810 150.945 ;
        RECT 60.340 150.915 61.340 150.945 ;
        RECT 56.770 150.660 57.000 150.805 ;
        RECT 57.970 150.660 58.200 150.805 ;
        RECT 58.945 150.660 59.205 150.735 ;
        RECT 59.905 150.660 60.135 150.805 ;
        RECT 61.545 150.660 61.775 150.805 ;
        RECT 61.930 150.690 62.230 150.945 ;
        RECT 62.985 150.945 64.540 151.115 ;
        RECT 67.030 151.050 68.935 151.115 ;
        RECT 69.695 151.115 69.985 152.190 ;
        RECT 70.190 152.160 70.420 152.305 ;
        RECT 71.390 152.160 71.620 152.305 ;
        RECT 72.335 152.160 72.655 152.205 ;
        RECT 73.325 152.160 73.555 152.305 ;
        RECT 74.965 152.160 75.195 152.305 ;
        RECT 70.190 151.990 75.195 152.160 ;
        RECT 70.190 151.845 70.420 151.990 ;
        RECT 71.390 151.845 71.620 151.990 ;
        RECT 72.335 151.945 72.655 151.990 ;
        RECT 73.325 151.845 73.555 151.990 ;
        RECT 74.965 151.845 75.195 151.990 ;
        RECT 70.580 151.705 71.230 151.735 ;
        RECT 72.365 151.705 72.625 151.780 ;
        RECT 73.760 151.705 74.760 151.735 ;
        RECT 70.560 151.535 74.780 151.705 ;
        RECT 70.580 151.505 71.230 151.535 ;
        RECT 72.365 151.460 72.625 151.535 ;
        RECT 73.300 151.375 73.470 151.535 ;
        RECT 73.760 151.505 74.760 151.535 ;
        RECT 70.580 151.115 71.230 151.145 ;
        RECT 67.030 150.945 68.940 151.050 ;
        RECT 56.770 150.490 61.775 150.660 ;
        RECT 56.770 150.345 57.000 150.490 ;
        RECT 57.970 150.345 58.200 150.490 ;
        RECT 58.945 150.415 59.205 150.490 ;
        RECT 59.905 150.345 60.135 150.490 ;
        RECT 61.545 150.345 61.775 150.490 ;
        RECT 57.140 150.235 57.400 150.280 ;
        RECT 57.140 150.205 57.810 150.235 ;
        RECT 60.340 150.205 61.340 150.235 ;
        RECT 57.140 150.035 61.360 150.205 ;
        RECT 57.140 150.005 57.810 150.035 ;
        RECT 60.340 150.005 61.340 150.035 ;
        RECT 57.140 149.960 57.400 150.005 ;
        RECT 57.160 149.615 57.810 149.645 ;
        RECT 60.340 149.615 61.340 149.645 ;
        RECT 61.935 149.615 62.225 150.690 ;
        RECT 56.275 149.550 57.830 149.615 ;
        RECT 49.560 149.190 49.860 149.445 ;
        RECT 50.450 149.415 51.100 149.445 ;
        RECT 53.630 149.415 54.630 149.445 ;
        RECT 49.565 148.115 49.855 149.190 ;
        RECT 50.060 149.160 50.290 149.305 ;
        RECT 51.260 149.160 51.490 149.305 ;
        RECT 53.195 149.235 53.425 149.305 ;
        RECT 53.130 149.160 53.425 149.235 ;
        RECT 54.835 149.160 55.065 149.305 ;
        RECT 50.060 148.990 55.065 149.160 ;
        RECT 50.060 148.845 50.290 148.990 ;
        RECT 51.260 148.845 51.490 148.990 ;
        RECT 53.130 148.915 53.425 148.990 ;
        RECT 53.195 148.845 53.425 148.915 ;
        RECT 54.835 148.845 55.065 148.990 ;
        RECT 50.450 148.705 51.100 148.735 ;
        RECT 52.235 148.705 52.495 148.780 ;
        RECT 53.630 148.705 54.630 148.735 ;
        RECT 50.430 148.535 52.495 148.705 ;
        RECT 53.610 148.535 54.650 148.705 ;
        RECT 50.450 148.505 51.100 148.535 ;
        RECT 52.235 148.460 52.495 148.535 ;
        RECT 53.630 148.505 54.630 148.535 ;
        RECT 54.045 148.145 54.215 148.505 ;
        RECT 50.450 148.115 51.100 148.145 ;
        RECT 53.630 148.115 54.630 148.145 ;
        RECT 36.640 147.490 41.645 147.660 ;
        RECT 36.640 147.345 36.870 147.490 ;
        RECT 37.840 147.345 38.070 147.490 ;
        RECT 39.775 147.345 40.005 147.490 ;
        RECT 40.550 147.415 40.810 147.490 ;
        RECT 41.415 147.345 41.645 147.490 ;
        RECT 37.030 147.205 37.680 147.235 ;
        RECT 38.815 147.205 39.075 147.280 ;
        RECT 40.210 147.205 41.210 147.235 ;
        RECT 37.010 147.035 39.075 147.205 ;
        RECT 40.190 147.035 41.230 147.205 ;
        RECT 37.030 147.005 37.680 147.035 ;
        RECT 38.815 146.960 39.075 147.035 ;
        RECT 40.210 147.005 41.210 147.035 ;
        RECT 40.625 146.645 40.795 147.005 ;
        RECT 37.030 146.615 37.680 146.645 ;
        RECT 40.210 146.615 41.210 146.645 ;
        RECT 36.145 146.550 37.700 146.615 ;
        RECT 36.140 146.445 37.700 146.550 ;
        RECT 40.190 146.445 41.230 146.615 ;
        RECT 36.140 146.190 36.440 146.445 ;
        RECT 37.030 146.415 37.680 146.445 ;
        RECT 40.210 146.415 41.210 146.445 ;
        RECT 36.145 145.115 36.435 146.190 ;
        RECT 36.640 146.160 36.870 146.305 ;
        RECT 37.840 146.160 38.070 146.305 ;
        RECT 39.775 146.160 40.005 146.305 ;
        RECT 40.970 146.160 41.230 146.235 ;
        RECT 41.415 146.160 41.645 146.305 ;
        RECT 36.640 145.990 41.645 146.160 ;
        RECT 36.640 145.845 36.870 145.990 ;
        RECT 37.840 145.845 38.070 145.990 ;
        RECT 39.775 145.845 40.005 145.990 ;
        RECT 40.970 145.915 41.230 145.990 ;
        RECT 41.415 145.845 41.645 145.990 ;
        RECT 37.030 145.705 37.680 145.735 ;
        RECT 38.815 145.705 39.075 145.780 ;
        RECT 40.210 145.705 41.210 145.735 ;
        RECT 37.010 145.535 41.230 145.705 ;
        RECT 37.030 145.505 37.680 145.535 ;
        RECT 38.815 145.460 39.075 145.535 ;
        RECT 40.210 145.505 41.210 145.535 ;
        RECT 37.030 145.115 37.680 145.145 ;
        RECT 40.210 145.115 41.210 145.145 ;
        RECT 41.805 145.115 42.095 147.690 ;
        RECT 42.855 146.615 43.145 147.945 ;
        RECT 43.740 147.915 44.390 147.945 ;
        RECT 46.920 147.915 47.920 147.945 ;
        RECT 43.350 147.660 43.580 147.805 ;
        RECT 44.550 147.660 44.780 147.805 ;
        RECT 46.485 147.660 46.715 147.805 ;
        RECT 47.260 147.660 47.520 147.735 ;
        RECT 48.125 147.660 48.355 147.805 ;
        RECT 48.510 147.690 48.810 148.050 ;
        RECT 49.565 147.945 51.120 148.115 ;
        RECT 53.610 147.945 54.650 148.115 ;
        RECT 55.225 148.050 55.515 149.445 ;
        RECT 56.270 149.445 57.830 149.550 ;
        RECT 60.320 149.445 62.225 149.615 ;
        RECT 62.985 149.615 63.275 150.945 ;
        RECT 63.870 150.915 64.520 150.945 ;
        RECT 67.050 150.915 68.050 150.945 ;
        RECT 63.480 150.660 63.710 150.805 ;
        RECT 64.680 150.660 64.910 150.805 ;
        RECT 65.655 150.660 65.915 150.735 ;
        RECT 66.615 150.660 66.845 150.805 ;
        RECT 68.255 150.660 68.485 150.805 ;
        RECT 68.640 150.690 68.940 150.945 ;
        RECT 69.695 150.945 71.250 151.115 ;
        RECT 73.255 151.055 73.515 151.375 ;
        RECT 73.760 151.115 74.760 151.145 ;
        RECT 75.355 151.115 75.645 152.445 ;
        RECT 76.400 152.445 77.960 152.550 ;
        RECT 80.450 152.445 82.355 152.615 ;
        RECT 83.115 153.660 83.405 153.945 ;
        RECT 84.000 153.915 84.650 153.945 ;
        RECT 87.180 153.915 88.180 153.945 ;
        RECT 83.610 153.660 83.840 153.805 ;
        RECT 84.810 153.660 85.040 153.805 ;
        RECT 86.745 153.660 86.975 153.805 ;
        RECT 88.385 153.660 88.615 153.805 ;
        RECT 88.770 153.690 89.070 153.945 ;
        RECT 89.825 153.945 91.380 154.115 ;
        RECT 93.870 154.050 95.775 154.115 ;
        RECT 96.535 154.115 96.825 154.325 ;
        RECT 97.420 154.115 98.070 154.145 ;
        RECT 100.600 154.115 101.600 154.145 ;
        RECT 102.195 154.115 102.485 154.325 ;
        RECT 93.870 153.945 95.780 154.050 ;
        RECT 83.115 153.490 88.615 153.660 ;
        RECT 83.115 152.615 83.405 153.490 ;
        RECT 83.610 153.345 83.840 153.490 ;
        RECT 84.810 153.345 85.040 153.490 ;
        RECT 86.745 153.345 86.975 153.490 ;
        RECT 88.385 153.345 88.615 153.490 ;
        RECT 84.000 153.205 84.650 153.235 ;
        RECT 87.180 153.205 88.180 153.235 ;
        RECT 83.980 153.035 88.200 153.205 ;
        RECT 84.000 153.005 84.650 153.035 ;
        RECT 87.180 153.005 88.180 153.035 ;
        RECT 84.000 152.615 84.650 152.645 ;
        RECT 87.180 152.615 88.180 152.645 ;
        RECT 88.775 152.615 89.065 153.690 ;
        RECT 83.115 152.550 84.670 152.615 ;
        RECT 76.400 152.190 76.700 152.445 ;
        RECT 77.290 152.415 77.940 152.445 ;
        RECT 80.470 152.415 81.470 152.445 ;
        RECT 73.740 151.050 75.645 151.115 ;
        RECT 76.405 151.115 76.695 152.190 ;
        RECT 76.900 152.160 77.130 152.305 ;
        RECT 78.100 152.160 78.330 152.305 ;
        RECT 79.045 152.160 79.365 152.205 ;
        RECT 80.035 152.160 80.265 152.305 ;
        RECT 81.675 152.160 81.905 152.305 ;
        RECT 76.900 151.990 81.905 152.160 ;
        RECT 76.900 151.845 77.130 151.990 ;
        RECT 78.100 151.845 78.330 151.990 ;
        RECT 79.045 151.945 79.365 151.990 ;
        RECT 80.035 151.845 80.265 151.990 ;
        RECT 81.675 151.845 81.905 151.990 ;
        RECT 77.290 151.705 77.940 151.735 ;
        RECT 79.075 151.705 79.335 151.780 ;
        RECT 80.390 151.735 80.650 151.780 ;
        RECT 80.390 151.705 81.470 151.735 ;
        RECT 77.270 151.535 81.490 151.705 ;
        RECT 77.290 151.505 77.940 151.535 ;
        RECT 79.075 151.460 79.335 151.535 ;
        RECT 80.390 151.505 81.470 151.535 ;
        RECT 80.390 151.460 80.650 151.505 ;
        RECT 77.290 151.115 77.940 151.145 ;
        RECT 80.470 151.115 81.470 151.145 ;
        RECT 82.065 151.115 82.355 152.445 ;
        RECT 83.110 152.445 84.670 152.550 ;
        RECT 87.160 152.445 89.065 152.615 ;
        RECT 89.825 152.615 90.115 153.945 ;
        RECT 90.710 153.915 91.360 153.945 ;
        RECT 93.890 153.915 94.890 153.945 ;
        RECT 90.320 153.660 90.550 153.805 ;
        RECT 90.690 153.660 90.950 153.735 ;
        RECT 91.520 153.660 91.750 153.805 ;
        RECT 93.455 153.660 93.685 153.805 ;
        RECT 95.095 153.660 95.325 153.805 ;
        RECT 95.480 153.690 95.780 153.945 ;
        RECT 96.535 153.945 98.090 154.115 ;
        RECT 100.580 154.050 102.485 154.115 ;
        RECT 100.580 153.945 102.490 154.050 ;
        RECT 90.320 153.490 95.325 153.660 ;
        RECT 90.320 153.345 90.550 153.490 ;
        RECT 90.690 153.415 90.950 153.490 ;
        RECT 91.520 153.345 91.750 153.490 ;
        RECT 93.455 153.345 93.685 153.490 ;
        RECT 95.095 153.345 95.325 153.490 ;
        RECT 94.650 153.235 94.910 153.280 ;
        RECT 90.710 153.205 91.360 153.235 ;
        RECT 93.890 153.205 94.910 153.235 ;
        RECT 90.690 153.035 94.910 153.205 ;
        RECT 90.710 153.005 91.360 153.035 ;
        RECT 93.890 153.005 94.910 153.035 ;
        RECT 94.650 152.960 94.910 153.005 ;
        RECT 90.710 152.615 91.360 152.645 ;
        RECT 93.890 152.615 94.890 152.645 ;
        RECT 95.485 152.615 95.775 153.690 ;
        RECT 89.825 152.550 91.380 152.615 ;
        RECT 83.110 152.190 83.410 152.445 ;
        RECT 84.000 152.415 84.650 152.445 ;
        RECT 87.180 152.415 88.180 152.445 ;
        RECT 73.740 150.945 75.650 151.050 ;
        RECT 63.480 150.490 68.485 150.660 ;
        RECT 63.480 150.345 63.710 150.490 ;
        RECT 64.680 150.345 64.910 150.490 ;
        RECT 65.655 150.415 65.915 150.490 ;
        RECT 66.615 150.345 66.845 150.490 ;
        RECT 68.255 150.345 68.485 150.490 ;
        RECT 67.390 150.235 67.650 150.280 ;
        RECT 63.870 150.205 64.520 150.235 ;
        RECT 67.050 150.205 68.050 150.235 ;
        RECT 63.850 150.035 68.070 150.205 ;
        RECT 63.870 150.005 64.520 150.035 ;
        RECT 67.050 150.005 68.050 150.035 ;
        RECT 67.390 149.960 67.650 150.005 ;
        RECT 63.870 149.615 64.520 149.645 ;
        RECT 67.050 149.615 68.050 149.645 ;
        RECT 68.645 149.615 68.935 150.690 ;
        RECT 62.985 149.550 64.540 149.615 ;
        RECT 56.270 149.190 56.570 149.445 ;
        RECT 57.160 149.415 57.810 149.445 ;
        RECT 60.340 149.415 61.340 149.445 ;
        RECT 56.275 148.115 56.565 149.190 ;
        RECT 56.770 149.160 57.000 149.305 ;
        RECT 57.970 149.160 58.200 149.305 ;
        RECT 59.905 149.235 60.135 149.305 ;
        RECT 59.840 149.160 60.135 149.235 ;
        RECT 61.545 149.160 61.775 149.305 ;
        RECT 56.770 148.990 61.775 149.160 ;
        RECT 56.770 148.845 57.000 148.990 ;
        RECT 57.970 148.845 58.200 148.990 ;
        RECT 59.840 148.915 60.135 148.990 ;
        RECT 59.905 148.845 60.135 148.915 ;
        RECT 61.545 148.845 61.775 148.990 ;
        RECT 57.160 148.705 57.810 148.735 ;
        RECT 58.945 148.705 59.205 148.780 ;
        RECT 60.340 148.705 61.340 148.735 ;
        RECT 57.140 148.535 59.205 148.705 ;
        RECT 60.320 148.535 61.360 148.705 ;
        RECT 57.160 148.505 57.810 148.535 ;
        RECT 58.945 148.460 59.205 148.535 ;
        RECT 60.340 148.505 61.340 148.535 ;
        RECT 60.755 148.145 60.925 148.505 ;
        RECT 57.160 148.115 57.810 148.145 ;
        RECT 60.340 148.115 61.340 148.145 ;
        RECT 43.350 147.490 48.355 147.660 ;
        RECT 43.350 147.345 43.580 147.490 ;
        RECT 44.550 147.345 44.780 147.490 ;
        RECT 46.485 147.345 46.715 147.490 ;
        RECT 47.260 147.415 47.520 147.490 ;
        RECT 48.125 147.345 48.355 147.490 ;
        RECT 43.740 147.205 44.390 147.235 ;
        RECT 45.525 147.205 45.785 147.280 ;
        RECT 46.920 147.205 47.920 147.235 ;
        RECT 43.720 147.035 45.785 147.205 ;
        RECT 46.900 147.035 47.940 147.205 ;
        RECT 43.740 147.005 44.390 147.035 ;
        RECT 45.525 146.960 45.785 147.035 ;
        RECT 46.920 147.005 47.920 147.035 ;
        RECT 47.335 146.645 47.505 147.005 ;
        RECT 43.740 146.615 44.390 146.645 ;
        RECT 46.920 146.615 47.920 146.645 ;
        RECT 42.855 146.550 44.410 146.615 ;
        RECT 42.850 146.445 44.410 146.550 ;
        RECT 46.900 146.445 47.940 146.615 ;
        RECT 42.850 146.190 43.150 146.445 ;
        RECT 43.740 146.415 44.390 146.445 ;
        RECT 46.920 146.415 47.920 146.445 ;
        RECT 36.145 144.945 37.700 145.115 ;
        RECT 40.190 145.050 42.095 145.115 ;
        RECT 42.855 145.115 43.145 146.190 ;
        RECT 43.350 146.160 43.580 146.305 ;
        RECT 44.550 146.160 44.780 146.305 ;
        RECT 46.485 146.160 46.715 146.305 ;
        RECT 47.680 146.160 47.940 146.235 ;
        RECT 48.125 146.160 48.355 146.305 ;
        RECT 43.350 145.990 48.355 146.160 ;
        RECT 43.350 145.845 43.580 145.990 ;
        RECT 44.550 145.845 44.780 145.990 ;
        RECT 46.485 145.845 46.715 145.990 ;
        RECT 47.680 145.915 47.940 145.990 ;
        RECT 48.125 145.845 48.355 145.990 ;
        RECT 43.740 145.705 44.390 145.735 ;
        RECT 45.525 145.705 45.785 145.780 ;
        RECT 46.920 145.705 47.920 145.735 ;
        RECT 43.720 145.535 47.940 145.705 ;
        RECT 43.740 145.505 44.390 145.535 ;
        RECT 45.525 145.460 45.785 145.535 ;
        RECT 46.920 145.505 47.920 145.535 ;
        RECT 43.740 145.115 44.390 145.145 ;
        RECT 46.920 145.115 47.920 145.145 ;
        RECT 48.515 145.115 48.805 147.690 ;
        RECT 49.565 146.615 49.855 147.945 ;
        RECT 50.450 147.915 51.100 147.945 ;
        RECT 53.630 147.915 54.630 147.945 ;
        RECT 50.060 147.660 50.290 147.805 ;
        RECT 51.260 147.660 51.490 147.805 ;
        RECT 53.195 147.660 53.425 147.805 ;
        RECT 53.970 147.660 54.230 147.735 ;
        RECT 54.835 147.660 55.065 147.805 ;
        RECT 55.220 147.690 55.520 148.050 ;
        RECT 56.275 147.945 57.830 148.115 ;
        RECT 60.320 147.945 61.360 148.115 ;
        RECT 61.935 148.050 62.225 149.445 ;
        RECT 62.980 149.445 64.540 149.550 ;
        RECT 67.030 149.445 68.935 149.615 ;
        RECT 69.695 149.615 69.985 150.945 ;
        RECT 70.580 150.915 71.230 150.945 ;
        RECT 73.760 150.915 74.760 150.945 ;
        RECT 70.190 150.660 70.420 150.805 ;
        RECT 71.390 150.660 71.620 150.805 ;
        RECT 72.365 150.660 72.625 150.735 ;
        RECT 73.325 150.660 73.555 150.805 ;
        RECT 74.965 150.660 75.195 150.805 ;
        RECT 75.350 150.690 75.650 150.945 ;
        RECT 76.405 150.945 77.960 151.115 ;
        RECT 80.450 151.050 82.355 151.115 ;
        RECT 83.115 151.115 83.405 152.190 ;
        RECT 83.610 152.160 83.840 152.305 ;
        RECT 84.810 152.160 85.040 152.305 ;
        RECT 85.755 152.160 86.075 152.205 ;
        RECT 86.745 152.160 86.975 152.305 ;
        RECT 88.385 152.160 88.615 152.305 ;
        RECT 83.610 151.990 88.615 152.160 ;
        RECT 83.610 151.845 83.840 151.990 ;
        RECT 84.810 151.845 85.040 151.990 ;
        RECT 85.755 151.945 86.075 151.990 ;
        RECT 86.745 151.845 86.975 151.990 ;
        RECT 88.385 151.845 88.615 151.990 ;
        RECT 84.000 151.705 84.650 151.735 ;
        RECT 85.785 151.705 86.045 151.780 ;
        RECT 87.180 151.705 88.180 151.735 ;
        RECT 83.980 151.535 88.200 151.705 ;
        RECT 84.000 151.505 84.650 151.535 ;
        RECT 85.785 151.460 86.045 151.535 ;
        RECT 86.720 151.375 86.890 151.535 ;
        RECT 87.180 151.505 88.180 151.535 ;
        RECT 84.000 151.115 84.650 151.145 ;
        RECT 80.450 150.945 82.360 151.050 ;
        RECT 70.190 150.490 75.195 150.660 ;
        RECT 70.190 150.345 70.420 150.490 ;
        RECT 71.390 150.345 71.620 150.490 ;
        RECT 72.365 150.415 72.625 150.490 ;
        RECT 73.325 150.345 73.555 150.490 ;
        RECT 74.965 150.345 75.195 150.490 ;
        RECT 70.560 150.235 70.820 150.280 ;
        RECT 70.560 150.205 71.230 150.235 ;
        RECT 73.760 150.205 74.760 150.235 ;
        RECT 70.560 150.035 74.780 150.205 ;
        RECT 70.560 150.005 71.230 150.035 ;
        RECT 73.760 150.005 74.760 150.035 ;
        RECT 70.560 149.960 70.820 150.005 ;
        RECT 70.580 149.615 71.230 149.645 ;
        RECT 73.760 149.615 74.760 149.645 ;
        RECT 75.355 149.615 75.645 150.690 ;
        RECT 69.695 149.550 71.250 149.615 ;
        RECT 62.980 149.190 63.280 149.445 ;
        RECT 63.870 149.415 64.520 149.445 ;
        RECT 67.050 149.415 68.050 149.445 ;
        RECT 62.985 148.115 63.275 149.190 ;
        RECT 63.480 149.160 63.710 149.305 ;
        RECT 64.680 149.160 64.910 149.305 ;
        RECT 66.615 149.235 66.845 149.305 ;
        RECT 66.550 149.160 66.845 149.235 ;
        RECT 68.255 149.160 68.485 149.305 ;
        RECT 63.480 148.990 68.485 149.160 ;
        RECT 63.480 148.845 63.710 148.990 ;
        RECT 64.680 148.845 64.910 148.990 ;
        RECT 66.550 148.915 66.845 148.990 ;
        RECT 66.615 148.845 66.845 148.915 ;
        RECT 68.255 148.845 68.485 148.990 ;
        RECT 63.870 148.705 64.520 148.735 ;
        RECT 65.655 148.705 65.915 148.780 ;
        RECT 67.050 148.705 68.050 148.735 ;
        RECT 63.850 148.535 65.915 148.705 ;
        RECT 67.030 148.535 68.070 148.705 ;
        RECT 63.870 148.505 64.520 148.535 ;
        RECT 65.655 148.460 65.915 148.535 ;
        RECT 67.050 148.505 68.050 148.535 ;
        RECT 67.465 148.145 67.635 148.505 ;
        RECT 63.870 148.115 64.520 148.145 ;
        RECT 67.050 148.115 68.050 148.145 ;
        RECT 50.060 147.490 55.065 147.660 ;
        RECT 50.060 147.345 50.290 147.490 ;
        RECT 51.260 147.345 51.490 147.490 ;
        RECT 53.195 147.345 53.425 147.490 ;
        RECT 53.970 147.415 54.230 147.490 ;
        RECT 54.835 147.345 55.065 147.490 ;
        RECT 50.450 147.205 51.100 147.235 ;
        RECT 52.235 147.205 52.495 147.280 ;
        RECT 53.630 147.205 54.630 147.235 ;
        RECT 50.430 147.035 52.495 147.205 ;
        RECT 53.610 147.035 54.650 147.205 ;
        RECT 50.450 147.005 51.100 147.035 ;
        RECT 52.235 146.960 52.495 147.035 ;
        RECT 53.630 147.005 54.630 147.035 ;
        RECT 54.045 146.645 54.215 147.005 ;
        RECT 50.450 146.615 51.100 146.645 ;
        RECT 53.630 146.615 54.630 146.645 ;
        RECT 49.565 146.550 51.120 146.615 ;
        RECT 49.560 146.445 51.120 146.550 ;
        RECT 53.610 146.445 54.650 146.615 ;
        RECT 49.560 146.190 49.860 146.445 ;
        RECT 50.450 146.415 51.100 146.445 ;
        RECT 53.630 146.415 54.630 146.445 ;
        RECT 40.190 144.945 42.100 145.050 ;
        RECT 36.145 143.615 36.435 144.945 ;
        RECT 37.030 144.915 37.680 144.945 ;
        RECT 40.210 144.915 41.210 144.945 ;
        RECT 36.640 144.660 36.870 144.805 ;
        RECT 37.840 144.660 38.070 144.805 ;
        RECT 39.775 144.735 40.005 144.805 ;
        RECT 39.710 144.660 40.005 144.735 ;
        RECT 41.415 144.660 41.645 144.805 ;
        RECT 41.800 144.690 42.100 144.945 ;
        RECT 42.855 144.945 44.410 145.115 ;
        RECT 46.900 145.050 48.805 145.115 ;
        RECT 49.565 145.115 49.855 146.190 ;
        RECT 50.060 146.160 50.290 146.305 ;
        RECT 51.260 146.160 51.490 146.305 ;
        RECT 53.195 146.160 53.425 146.305 ;
        RECT 54.390 146.160 54.650 146.235 ;
        RECT 54.835 146.160 55.065 146.305 ;
        RECT 50.060 145.990 55.065 146.160 ;
        RECT 50.060 145.845 50.290 145.990 ;
        RECT 51.260 145.845 51.490 145.990 ;
        RECT 53.195 145.845 53.425 145.990 ;
        RECT 54.390 145.915 54.650 145.990 ;
        RECT 54.835 145.845 55.065 145.990 ;
        RECT 50.450 145.705 51.100 145.735 ;
        RECT 52.235 145.705 52.495 145.780 ;
        RECT 53.630 145.705 54.630 145.735 ;
        RECT 50.430 145.535 54.650 145.705 ;
        RECT 50.450 145.505 51.100 145.535 ;
        RECT 52.235 145.460 52.495 145.535 ;
        RECT 53.630 145.505 54.630 145.535 ;
        RECT 50.450 145.115 51.100 145.145 ;
        RECT 53.630 145.115 54.630 145.145 ;
        RECT 55.225 145.115 55.515 147.690 ;
        RECT 56.275 146.615 56.565 147.945 ;
        RECT 57.160 147.915 57.810 147.945 ;
        RECT 60.340 147.915 61.340 147.945 ;
        RECT 56.770 147.660 57.000 147.805 ;
        RECT 57.970 147.660 58.200 147.805 ;
        RECT 59.905 147.660 60.135 147.805 ;
        RECT 60.680 147.660 60.940 147.735 ;
        RECT 61.545 147.660 61.775 147.805 ;
        RECT 61.930 147.690 62.230 148.050 ;
        RECT 62.985 147.945 64.540 148.115 ;
        RECT 67.030 147.945 68.070 148.115 ;
        RECT 68.645 148.050 68.935 149.445 ;
        RECT 69.690 149.445 71.250 149.550 ;
        RECT 73.740 149.445 75.645 149.615 ;
        RECT 76.405 149.615 76.695 150.945 ;
        RECT 77.290 150.915 77.940 150.945 ;
        RECT 80.470 150.915 81.470 150.945 ;
        RECT 76.900 150.660 77.130 150.805 ;
        RECT 78.100 150.660 78.330 150.805 ;
        RECT 79.075 150.660 79.335 150.735 ;
        RECT 80.035 150.660 80.265 150.805 ;
        RECT 81.675 150.660 81.905 150.805 ;
        RECT 82.060 150.690 82.360 150.945 ;
        RECT 83.115 150.945 84.670 151.115 ;
        RECT 86.675 151.055 86.935 151.375 ;
        RECT 87.180 151.115 88.180 151.145 ;
        RECT 88.775 151.115 89.065 152.445 ;
        RECT 89.820 152.445 91.380 152.550 ;
        RECT 93.870 152.445 95.775 152.615 ;
        RECT 96.535 153.660 96.825 153.945 ;
        RECT 97.420 153.915 98.070 153.945 ;
        RECT 100.600 153.915 101.600 153.945 ;
        RECT 97.030 153.660 97.260 153.805 ;
        RECT 98.230 153.660 98.460 153.805 ;
        RECT 100.165 153.660 100.395 153.805 ;
        RECT 101.805 153.660 102.035 153.805 ;
        RECT 102.190 153.690 102.490 153.945 ;
        RECT 96.535 153.490 102.035 153.660 ;
        RECT 96.535 152.615 96.825 153.490 ;
        RECT 97.030 153.345 97.260 153.490 ;
        RECT 98.230 153.345 98.460 153.490 ;
        RECT 100.165 153.345 100.395 153.490 ;
        RECT 101.805 153.345 102.035 153.490 ;
        RECT 97.420 153.205 98.070 153.235 ;
        RECT 100.600 153.205 101.600 153.235 ;
        RECT 97.400 153.035 101.620 153.205 ;
        RECT 97.420 153.005 98.070 153.035 ;
        RECT 100.600 153.005 101.600 153.035 ;
        RECT 97.420 152.615 98.070 152.645 ;
        RECT 100.600 152.615 101.600 152.645 ;
        RECT 102.195 152.615 102.485 153.690 ;
        RECT 96.535 152.550 98.090 152.615 ;
        RECT 89.820 152.190 90.120 152.445 ;
        RECT 90.710 152.415 91.360 152.445 ;
        RECT 93.890 152.415 94.890 152.445 ;
        RECT 87.160 151.050 89.065 151.115 ;
        RECT 89.825 151.115 90.115 152.190 ;
        RECT 90.320 152.160 90.550 152.305 ;
        RECT 91.520 152.160 91.750 152.305 ;
        RECT 92.465 152.160 92.785 152.205 ;
        RECT 93.455 152.160 93.685 152.305 ;
        RECT 95.095 152.160 95.325 152.305 ;
        RECT 90.320 151.990 95.325 152.160 ;
        RECT 90.320 151.845 90.550 151.990 ;
        RECT 91.520 151.845 91.750 151.990 ;
        RECT 92.465 151.945 92.785 151.990 ;
        RECT 93.455 151.845 93.685 151.990 ;
        RECT 95.095 151.845 95.325 151.990 ;
        RECT 90.710 151.705 91.360 151.735 ;
        RECT 92.495 151.705 92.755 151.780 ;
        RECT 93.810 151.735 94.070 151.780 ;
        RECT 93.810 151.705 94.890 151.735 ;
        RECT 90.690 151.535 94.910 151.705 ;
        RECT 90.710 151.505 91.360 151.535 ;
        RECT 92.495 151.460 92.755 151.535 ;
        RECT 93.810 151.505 94.890 151.535 ;
        RECT 93.810 151.460 94.070 151.505 ;
        RECT 90.710 151.115 91.360 151.145 ;
        RECT 93.890 151.115 94.890 151.145 ;
        RECT 95.485 151.115 95.775 152.445 ;
        RECT 96.530 152.445 98.090 152.550 ;
        RECT 100.580 152.445 102.485 152.615 ;
        RECT 96.530 152.190 96.830 152.445 ;
        RECT 97.420 152.415 98.070 152.445 ;
        RECT 100.600 152.415 101.600 152.445 ;
        RECT 87.160 150.945 89.070 151.050 ;
        RECT 76.900 150.490 81.905 150.660 ;
        RECT 76.900 150.345 77.130 150.490 ;
        RECT 78.100 150.345 78.330 150.490 ;
        RECT 79.075 150.415 79.335 150.490 ;
        RECT 80.035 150.345 80.265 150.490 ;
        RECT 81.675 150.345 81.905 150.490 ;
        RECT 80.810 150.235 81.070 150.280 ;
        RECT 77.290 150.205 77.940 150.235 ;
        RECT 80.470 150.205 81.470 150.235 ;
        RECT 77.270 150.035 81.490 150.205 ;
        RECT 77.290 150.005 77.940 150.035 ;
        RECT 80.470 150.005 81.470 150.035 ;
        RECT 80.810 149.960 81.070 150.005 ;
        RECT 77.290 149.615 77.940 149.645 ;
        RECT 80.470 149.615 81.470 149.645 ;
        RECT 82.065 149.615 82.355 150.690 ;
        RECT 76.405 149.550 77.960 149.615 ;
        RECT 69.690 149.190 69.990 149.445 ;
        RECT 70.580 149.415 71.230 149.445 ;
        RECT 73.760 149.415 74.760 149.445 ;
        RECT 69.695 148.115 69.985 149.190 ;
        RECT 70.190 149.160 70.420 149.305 ;
        RECT 71.390 149.160 71.620 149.305 ;
        RECT 73.325 149.235 73.555 149.305 ;
        RECT 73.260 149.160 73.555 149.235 ;
        RECT 74.965 149.160 75.195 149.305 ;
        RECT 70.190 148.990 75.195 149.160 ;
        RECT 70.190 148.845 70.420 148.990 ;
        RECT 71.390 148.845 71.620 148.990 ;
        RECT 73.260 148.915 73.555 148.990 ;
        RECT 73.325 148.845 73.555 148.915 ;
        RECT 74.965 148.845 75.195 148.990 ;
        RECT 70.580 148.705 71.230 148.735 ;
        RECT 72.365 148.705 72.625 148.780 ;
        RECT 73.760 148.705 74.760 148.735 ;
        RECT 70.560 148.535 72.625 148.705 ;
        RECT 73.740 148.535 74.780 148.705 ;
        RECT 70.580 148.505 71.230 148.535 ;
        RECT 72.365 148.460 72.625 148.535 ;
        RECT 73.760 148.505 74.760 148.535 ;
        RECT 74.175 148.145 74.345 148.505 ;
        RECT 70.580 148.115 71.230 148.145 ;
        RECT 73.760 148.115 74.760 148.145 ;
        RECT 56.770 147.490 61.775 147.660 ;
        RECT 56.770 147.345 57.000 147.490 ;
        RECT 57.970 147.345 58.200 147.490 ;
        RECT 59.905 147.345 60.135 147.490 ;
        RECT 60.680 147.415 60.940 147.490 ;
        RECT 61.545 147.345 61.775 147.490 ;
        RECT 57.160 147.205 57.810 147.235 ;
        RECT 58.945 147.205 59.205 147.280 ;
        RECT 60.340 147.205 61.340 147.235 ;
        RECT 57.140 147.035 59.205 147.205 ;
        RECT 60.320 147.035 61.360 147.205 ;
        RECT 57.160 147.005 57.810 147.035 ;
        RECT 58.945 146.960 59.205 147.035 ;
        RECT 60.340 147.005 61.340 147.035 ;
        RECT 60.755 146.645 60.925 147.005 ;
        RECT 57.160 146.615 57.810 146.645 ;
        RECT 60.340 146.615 61.340 146.645 ;
        RECT 56.275 146.550 57.830 146.615 ;
        RECT 56.270 146.445 57.830 146.550 ;
        RECT 60.320 146.445 61.360 146.615 ;
        RECT 56.270 146.190 56.570 146.445 ;
        RECT 57.160 146.415 57.810 146.445 ;
        RECT 60.340 146.415 61.340 146.445 ;
        RECT 46.900 144.945 48.810 145.050 ;
        RECT 36.640 144.490 41.645 144.660 ;
        RECT 36.640 144.345 36.870 144.490 ;
        RECT 37.840 144.345 38.070 144.490 ;
        RECT 39.710 144.415 40.005 144.490 ;
        RECT 39.775 144.345 40.005 144.415 ;
        RECT 41.415 144.345 41.645 144.490 ;
        RECT 37.030 144.205 37.680 144.235 ;
        RECT 38.815 144.205 39.075 144.280 ;
        RECT 40.210 144.205 41.210 144.235 ;
        RECT 37.010 144.035 39.075 144.205 ;
        RECT 40.190 144.035 41.230 144.205 ;
        RECT 37.030 144.005 37.680 144.035 ;
        RECT 38.815 143.960 39.075 144.035 ;
        RECT 40.210 144.005 41.210 144.035 ;
        RECT 40.625 143.645 40.795 144.005 ;
        RECT 37.030 143.615 37.680 143.645 ;
        RECT 40.210 143.615 41.210 143.645 ;
        RECT 36.145 143.550 37.700 143.615 ;
        RECT 36.140 143.445 37.700 143.550 ;
        RECT 40.190 143.445 41.230 143.615 ;
        RECT 36.140 143.190 36.440 143.445 ;
        RECT 37.030 143.415 37.680 143.445 ;
        RECT 40.210 143.415 41.210 143.445 ;
        RECT 36.145 142.115 36.435 143.190 ;
        RECT 36.640 143.160 36.870 143.305 ;
        RECT 37.840 143.160 38.070 143.305 ;
        RECT 39.775 143.235 40.005 143.305 ;
        RECT 39.775 143.160 40.390 143.235 ;
        RECT 41.415 143.160 41.645 143.305 ;
        RECT 36.640 142.990 41.645 143.160 ;
        RECT 36.640 142.845 36.870 142.990 ;
        RECT 37.840 142.845 38.070 142.990 ;
        RECT 39.775 142.915 40.390 142.990 ;
        RECT 39.775 142.845 40.005 142.915 ;
        RECT 41.415 142.845 41.645 142.990 ;
        RECT 37.030 142.705 37.680 142.735 ;
        RECT 38.815 142.705 39.075 142.780 ;
        RECT 40.210 142.705 41.210 142.735 ;
        RECT 37.010 142.535 39.075 142.705 ;
        RECT 40.190 142.535 41.230 142.705 ;
        RECT 37.030 142.505 37.680 142.535 ;
        RECT 38.815 142.460 39.075 142.535 ;
        RECT 40.210 142.505 41.210 142.535 ;
        RECT 40.625 142.145 40.795 142.505 ;
        RECT 37.030 142.115 37.680 142.145 ;
        RECT 40.210 142.115 41.210 142.145 ;
        RECT 36.145 141.945 37.700 142.115 ;
        RECT 40.190 141.945 41.230 142.115 ;
        RECT 41.805 142.050 42.095 144.690 ;
        RECT 42.855 143.615 43.145 144.945 ;
        RECT 43.740 144.915 44.390 144.945 ;
        RECT 46.920 144.915 47.920 144.945 ;
        RECT 43.350 144.660 43.580 144.805 ;
        RECT 44.550 144.660 44.780 144.805 ;
        RECT 46.485 144.735 46.715 144.805 ;
        RECT 46.420 144.660 46.715 144.735 ;
        RECT 48.125 144.660 48.355 144.805 ;
        RECT 48.510 144.690 48.810 144.945 ;
        RECT 49.565 144.945 51.120 145.115 ;
        RECT 53.610 145.050 55.515 145.115 ;
        RECT 56.275 145.115 56.565 146.190 ;
        RECT 56.770 146.160 57.000 146.305 ;
        RECT 57.970 146.160 58.200 146.305 ;
        RECT 59.905 146.160 60.135 146.305 ;
        RECT 61.100 146.160 61.360 146.235 ;
        RECT 61.545 146.160 61.775 146.305 ;
        RECT 56.770 145.990 61.775 146.160 ;
        RECT 56.770 145.845 57.000 145.990 ;
        RECT 57.970 145.845 58.200 145.990 ;
        RECT 59.905 145.845 60.135 145.990 ;
        RECT 61.100 145.915 61.360 145.990 ;
        RECT 61.545 145.845 61.775 145.990 ;
        RECT 57.160 145.705 57.810 145.735 ;
        RECT 58.945 145.705 59.205 145.780 ;
        RECT 60.340 145.705 61.340 145.735 ;
        RECT 57.140 145.535 61.360 145.705 ;
        RECT 57.160 145.505 57.810 145.535 ;
        RECT 58.945 145.460 59.205 145.535 ;
        RECT 60.340 145.505 61.340 145.535 ;
        RECT 57.160 145.115 57.810 145.145 ;
        RECT 60.340 145.115 61.340 145.145 ;
        RECT 61.935 145.115 62.225 147.690 ;
        RECT 62.985 146.615 63.275 147.945 ;
        RECT 63.870 147.915 64.520 147.945 ;
        RECT 67.050 147.915 68.050 147.945 ;
        RECT 63.480 147.660 63.710 147.805 ;
        RECT 64.680 147.660 64.910 147.805 ;
        RECT 66.615 147.660 66.845 147.805 ;
        RECT 67.390 147.660 67.650 147.735 ;
        RECT 68.255 147.660 68.485 147.805 ;
        RECT 68.640 147.690 68.940 148.050 ;
        RECT 69.695 147.945 71.250 148.115 ;
        RECT 73.740 147.945 74.780 148.115 ;
        RECT 75.355 148.050 75.645 149.445 ;
        RECT 76.400 149.445 77.960 149.550 ;
        RECT 80.450 149.445 82.355 149.615 ;
        RECT 83.115 149.615 83.405 150.945 ;
        RECT 84.000 150.915 84.650 150.945 ;
        RECT 87.180 150.915 88.180 150.945 ;
        RECT 83.610 150.660 83.840 150.805 ;
        RECT 84.810 150.660 85.040 150.805 ;
        RECT 85.785 150.660 86.045 150.735 ;
        RECT 86.745 150.660 86.975 150.805 ;
        RECT 88.385 150.660 88.615 150.805 ;
        RECT 88.770 150.690 89.070 150.945 ;
        RECT 89.825 150.945 91.380 151.115 ;
        RECT 93.870 151.050 95.775 151.115 ;
        RECT 96.535 151.115 96.825 152.190 ;
        RECT 97.030 152.160 97.260 152.305 ;
        RECT 98.230 152.160 98.460 152.305 ;
        RECT 99.175 152.160 99.495 152.205 ;
        RECT 100.165 152.160 100.395 152.305 ;
        RECT 101.805 152.160 102.035 152.305 ;
        RECT 97.030 151.990 102.035 152.160 ;
        RECT 97.030 151.845 97.260 151.990 ;
        RECT 98.230 151.845 98.460 151.990 ;
        RECT 99.175 151.945 99.495 151.990 ;
        RECT 100.165 151.845 100.395 151.990 ;
        RECT 101.805 151.845 102.035 151.990 ;
        RECT 97.420 151.705 98.070 151.735 ;
        RECT 99.205 151.705 99.465 151.780 ;
        RECT 100.600 151.705 101.600 151.735 ;
        RECT 97.400 151.535 101.620 151.705 ;
        RECT 97.420 151.505 98.070 151.535 ;
        RECT 99.205 151.460 99.465 151.535 ;
        RECT 100.140 151.375 100.310 151.535 ;
        RECT 100.600 151.505 101.600 151.535 ;
        RECT 97.420 151.115 98.070 151.145 ;
        RECT 93.870 150.945 95.780 151.050 ;
        RECT 83.610 150.490 88.615 150.660 ;
        RECT 83.610 150.345 83.840 150.490 ;
        RECT 84.810 150.345 85.040 150.490 ;
        RECT 85.785 150.415 86.045 150.490 ;
        RECT 86.745 150.345 86.975 150.490 ;
        RECT 88.385 150.345 88.615 150.490 ;
        RECT 83.980 150.235 84.240 150.280 ;
        RECT 83.980 150.205 84.650 150.235 ;
        RECT 87.180 150.205 88.180 150.235 ;
        RECT 83.980 150.035 88.200 150.205 ;
        RECT 83.980 150.005 84.650 150.035 ;
        RECT 87.180 150.005 88.180 150.035 ;
        RECT 83.980 149.960 84.240 150.005 ;
        RECT 84.000 149.615 84.650 149.645 ;
        RECT 87.180 149.615 88.180 149.645 ;
        RECT 88.775 149.615 89.065 150.690 ;
        RECT 83.115 149.550 84.670 149.615 ;
        RECT 76.400 149.190 76.700 149.445 ;
        RECT 77.290 149.415 77.940 149.445 ;
        RECT 80.470 149.415 81.470 149.445 ;
        RECT 76.405 148.115 76.695 149.190 ;
        RECT 76.900 149.160 77.130 149.305 ;
        RECT 78.100 149.160 78.330 149.305 ;
        RECT 80.035 149.235 80.265 149.305 ;
        RECT 79.970 149.160 80.265 149.235 ;
        RECT 81.675 149.160 81.905 149.305 ;
        RECT 76.900 148.990 81.905 149.160 ;
        RECT 76.900 148.845 77.130 148.990 ;
        RECT 78.100 148.845 78.330 148.990 ;
        RECT 79.970 148.915 80.265 148.990 ;
        RECT 80.035 148.845 80.265 148.915 ;
        RECT 81.675 148.845 81.905 148.990 ;
        RECT 77.290 148.705 77.940 148.735 ;
        RECT 79.075 148.705 79.335 148.780 ;
        RECT 80.470 148.705 81.470 148.735 ;
        RECT 77.270 148.535 79.335 148.705 ;
        RECT 80.450 148.535 81.490 148.705 ;
        RECT 77.290 148.505 77.940 148.535 ;
        RECT 79.075 148.460 79.335 148.535 ;
        RECT 80.470 148.505 81.470 148.535 ;
        RECT 80.885 148.145 81.055 148.505 ;
        RECT 77.290 148.115 77.940 148.145 ;
        RECT 80.470 148.115 81.470 148.145 ;
        RECT 63.480 147.490 68.485 147.660 ;
        RECT 63.480 147.345 63.710 147.490 ;
        RECT 64.680 147.345 64.910 147.490 ;
        RECT 66.615 147.345 66.845 147.490 ;
        RECT 67.390 147.415 67.650 147.490 ;
        RECT 68.255 147.345 68.485 147.490 ;
        RECT 63.870 147.205 64.520 147.235 ;
        RECT 65.655 147.205 65.915 147.280 ;
        RECT 67.050 147.205 68.050 147.235 ;
        RECT 63.850 147.035 65.915 147.205 ;
        RECT 67.030 147.035 68.070 147.205 ;
        RECT 63.870 147.005 64.520 147.035 ;
        RECT 65.655 146.960 65.915 147.035 ;
        RECT 67.050 147.005 68.050 147.035 ;
        RECT 67.465 146.645 67.635 147.005 ;
        RECT 63.870 146.615 64.520 146.645 ;
        RECT 67.050 146.615 68.050 146.645 ;
        RECT 62.985 146.550 64.540 146.615 ;
        RECT 62.980 146.445 64.540 146.550 ;
        RECT 67.030 146.445 68.070 146.615 ;
        RECT 62.980 146.190 63.280 146.445 ;
        RECT 63.870 146.415 64.520 146.445 ;
        RECT 67.050 146.415 68.050 146.445 ;
        RECT 53.610 144.945 55.520 145.050 ;
        RECT 43.350 144.490 48.355 144.660 ;
        RECT 43.350 144.345 43.580 144.490 ;
        RECT 44.550 144.345 44.780 144.490 ;
        RECT 46.420 144.415 46.715 144.490 ;
        RECT 46.485 144.345 46.715 144.415 ;
        RECT 48.125 144.345 48.355 144.490 ;
        RECT 43.740 144.205 44.390 144.235 ;
        RECT 45.525 144.205 45.785 144.280 ;
        RECT 46.920 144.205 47.920 144.235 ;
        RECT 43.720 144.035 45.785 144.205 ;
        RECT 46.900 144.035 47.940 144.205 ;
        RECT 43.740 144.005 44.390 144.035 ;
        RECT 45.525 143.960 45.785 144.035 ;
        RECT 46.920 144.005 47.920 144.035 ;
        RECT 47.335 143.645 47.505 144.005 ;
        RECT 43.740 143.615 44.390 143.645 ;
        RECT 46.920 143.615 47.920 143.645 ;
        RECT 42.855 143.550 44.410 143.615 ;
        RECT 42.850 143.445 44.410 143.550 ;
        RECT 46.900 143.445 47.940 143.615 ;
        RECT 42.850 143.190 43.150 143.445 ;
        RECT 43.740 143.415 44.390 143.445 ;
        RECT 46.920 143.415 47.920 143.445 ;
        RECT 42.855 142.115 43.145 143.190 ;
        RECT 43.350 143.160 43.580 143.305 ;
        RECT 44.550 143.160 44.780 143.305 ;
        RECT 46.485 143.235 46.715 143.305 ;
        RECT 46.485 143.160 47.100 143.235 ;
        RECT 48.125 143.160 48.355 143.305 ;
        RECT 43.350 142.990 48.355 143.160 ;
        RECT 43.350 142.845 43.580 142.990 ;
        RECT 44.550 142.845 44.780 142.990 ;
        RECT 46.485 142.915 47.100 142.990 ;
        RECT 46.485 142.845 46.715 142.915 ;
        RECT 48.125 142.845 48.355 142.990 ;
        RECT 43.740 142.705 44.390 142.735 ;
        RECT 45.525 142.705 45.785 142.780 ;
        RECT 46.920 142.705 47.920 142.735 ;
        RECT 43.720 142.535 45.785 142.705 ;
        RECT 46.900 142.535 47.940 142.705 ;
        RECT 43.740 142.505 44.390 142.535 ;
        RECT 45.525 142.460 45.785 142.535 ;
        RECT 46.920 142.505 47.920 142.535 ;
        RECT 47.335 142.145 47.505 142.505 ;
        RECT 43.740 142.115 44.390 142.145 ;
        RECT 46.920 142.115 47.920 142.145 ;
        RECT 36.145 140.825 36.435 141.945 ;
        RECT 37.030 141.915 37.680 141.945 ;
        RECT 40.210 141.915 41.210 141.945 ;
        RECT 36.640 141.660 36.870 141.805 ;
        RECT 37.840 141.660 38.070 141.805 ;
        RECT 39.775 141.660 40.005 141.805 ;
        RECT 40.970 141.660 41.230 141.735 ;
        RECT 41.415 141.660 41.645 141.805 ;
        RECT 41.800 141.690 42.100 142.050 ;
        RECT 42.855 141.945 44.410 142.115 ;
        RECT 46.900 141.945 47.940 142.115 ;
        RECT 48.515 142.050 48.805 144.690 ;
        RECT 49.565 143.615 49.855 144.945 ;
        RECT 50.450 144.915 51.100 144.945 ;
        RECT 53.630 144.915 54.630 144.945 ;
        RECT 50.060 144.660 50.290 144.805 ;
        RECT 51.260 144.660 51.490 144.805 ;
        RECT 53.195 144.735 53.425 144.805 ;
        RECT 53.130 144.660 53.425 144.735 ;
        RECT 54.835 144.660 55.065 144.805 ;
        RECT 55.220 144.690 55.520 144.945 ;
        RECT 56.275 144.945 57.830 145.115 ;
        RECT 60.320 145.050 62.225 145.115 ;
        RECT 62.985 145.115 63.275 146.190 ;
        RECT 63.480 146.160 63.710 146.305 ;
        RECT 64.680 146.160 64.910 146.305 ;
        RECT 66.615 146.160 66.845 146.305 ;
        RECT 67.810 146.160 68.070 146.235 ;
        RECT 68.255 146.160 68.485 146.305 ;
        RECT 63.480 145.990 68.485 146.160 ;
        RECT 63.480 145.845 63.710 145.990 ;
        RECT 64.680 145.845 64.910 145.990 ;
        RECT 66.615 145.845 66.845 145.990 ;
        RECT 67.810 145.915 68.070 145.990 ;
        RECT 68.255 145.845 68.485 145.990 ;
        RECT 63.870 145.705 64.520 145.735 ;
        RECT 65.655 145.705 65.915 145.780 ;
        RECT 67.050 145.705 68.050 145.735 ;
        RECT 63.850 145.535 68.070 145.705 ;
        RECT 63.870 145.505 64.520 145.535 ;
        RECT 65.655 145.460 65.915 145.535 ;
        RECT 67.050 145.505 68.050 145.535 ;
        RECT 63.870 145.115 64.520 145.145 ;
        RECT 67.050 145.115 68.050 145.145 ;
        RECT 68.645 145.115 68.935 147.690 ;
        RECT 69.695 146.615 69.985 147.945 ;
        RECT 70.580 147.915 71.230 147.945 ;
        RECT 73.760 147.915 74.760 147.945 ;
        RECT 70.190 147.660 70.420 147.805 ;
        RECT 71.390 147.660 71.620 147.805 ;
        RECT 73.325 147.660 73.555 147.805 ;
        RECT 74.100 147.660 74.360 147.735 ;
        RECT 74.965 147.660 75.195 147.805 ;
        RECT 75.350 147.690 75.650 148.050 ;
        RECT 76.405 147.945 77.960 148.115 ;
        RECT 80.450 147.945 81.490 148.115 ;
        RECT 82.065 148.050 82.355 149.445 ;
        RECT 83.110 149.445 84.670 149.550 ;
        RECT 87.160 149.445 89.065 149.615 ;
        RECT 89.825 149.615 90.115 150.945 ;
        RECT 90.710 150.915 91.360 150.945 ;
        RECT 93.890 150.915 94.890 150.945 ;
        RECT 90.320 150.660 90.550 150.805 ;
        RECT 91.520 150.660 91.750 150.805 ;
        RECT 92.495 150.660 92.755 150.735 ;
        RECT 93.455 150.660 93.685 150.805 ;
        RECT 95.095 150.660 95.325 150.805 ;
        RECT 95.480 150.690 95.780 150.945 ;
        RECT 96.535 150.945 98.090 151.115 ;
        RECT 100.095 151.055 100.355 151.375 ;
        RECT 100.600 151.115 101.600 151.145 ;
        RECT 102.195 151.115 102.485 152.445 ;
        RECT 100.580 151.050 102.485 151.115 ;
        RECT 100.580 150.945 102.490 151.050 ;
        RECT 90.320 150.490 95.325 150.660 ;
        RECT 90.320 150.345 90.550 150.490 ;
        RECT 91.520 150.345 91.750 150.490 ;
        RECT 92.495 150.415 92.755 150.490 ;
        RECT 93.455 150.345 93.685 150.490 ;
        RECT 95.095 150.345 95.325 150.490 ;
        RECT 94.230 150.235 94.490 150.280 ;
        RECT 90.710 150.205 91.360 150.235 ;
        RECT 93.890 150.205 94.890 150.235 ;
        RECT 90.690 150.035 94.910 150.205 ;
        RECT 90.710 150.005 91.360 150.035 ;
        RECT 93.890 150.005 94.890 150.035 ;
        RECT 94.230 149.960 94.490 150.005 ;
        RECT 90.710 149.615 91.360 149.645 ;
        RECT 93.890 149.615 94.890 149.645 ;
        RECT 95.485 149.615 95.775 150.690 ;
        RECT 89.825 149.550 91.380 149.615 ;
        RECT 83.110 149.190 83.410 149.445 ;
        RECT 84.000 149.415 84.650 149.445 ;
        RECT 87.180 149.415 88.180 149.445 ;
        RECT 83.115 148.115 83.405 149.190 ;
        RECT 83.610 149.160 83.840 149.305 ;
        RECT 84.810 149.160 85.040 149.305 ;
        RECT 86.745 149.235 86.975 149.305 ;
        RECT 86.680 149.160 86.975 149.235 ;
        RECT 88.385 149.160 88.615 149.305 ;
        RECT 83.610 148.990 88.615 149.160 ;
        RECT 83.610 148.845 83.840 148.990 ;
        RECT 84.810 148.845 85.040 148.990 ;
        RECT 86.680 148.915 86.975 148.990 ;
        RECT 86.745 148.845 86.975 148.915 ;
        RECT 88.385 148.845 88.615 148.990 ;
        RECT 84.000 148.705 84.650 148.735 ;
        RECT 85.785 148.705 86.045 148.780 ;
        RECT 87.180 148.705 88.180 148.735 ;
        RECT 83.980 148.535 86.045 148.705 ;
        RECT 87.160 148.535 88.200 148.705 ;
        RECT 84.000 148.505 84.650 148.535 ;
        RECT 85.785 148.460 86.045 148.535 ;
        RECT 87.180 148.505 88.180 148.535 ;
        RECT 87.595 148.145 87.765 148.505 ;
        RECT 84.000 148.115 84.650 148.145 ;
        RECT 87.180 148.115 88.180 148.145 ;
        RECT 70.190 147.490 75.195 147.660 ;
        RECT 70.190 147.345 70.420 147.490 ;
        RECT 71.390 147.345 71.620 147.490 ;
        RECT 73.325 147.345 73.555 147.490 ;
        RECT 74.100 147.415 74.360 147.490 ;
        RECT 74.965 147.345 75.195 147.490 ;
        RECT 70.580 147.205 71.230 147.235 ;
        RECT 72.365 147.205 72.625 147.280 ;
        RECT 73.760 147.205 74.760 147.235 ;
        RECT 70.560 147.035 72.625 147.205 ;
        RECT 73.740 147.035 74.780 147.205 ;
        RECT 70.580 147.005 71.230 147.035 ;
        RECT 72.365 146.960 72.625 147.035 ;
        RECT 73.760 147.005 74.760 147.035 ;
        RECT 74.175 146.645 74.345 147.005 ;
        RECT 70.580 146.615 71.230 146.645 ;
        RECT 73.760 146.615 74.760 146.645 ;
        RECT 69.695 146.550 71.250 146.615 ;
        RECT 69.690 146.445 71.250 146.550 ;
        RECT 73.740 146.445 74.780 146.615 ;
        RECT 69.690 146.190 69.990 146.445 ;
        RECT 70.580 146.415 71.230 146.445 ;
        RECT 73.760 146.415 74.760 146.445 ;
        RECT 60.320 144.945 62.230 145.050 ;
        RECT 50.060 144.490 55.065 144.660 ;
        RECT 50.060 144.345 50.290 144.490 ;
        RECT 51.260 144.345 51.490 144.490 ;
        RECT 53.130 144.415 53.425 144.490 ;
        RECT 53.195 144.345 53.425 144.415 ;
        RECT 54.835 144.345 55.065 144.490 ;
        RECT 50.450 144.205 51.100 144.235 ;
        RECT 52.235 144.205 52.495 144.280 ;
        RECT 53.630 144.205 54.630 144.235 ;
        RECT 50.430 144.035 52.495 144.205 ;
        RECT 53.610 144.035 54.650 144.205 ;
        RECT 50.450 144.005 51.100 144.035 ;
        RECT 52.235 143.960 52.495 144.035 ;
        RECT 53.630 144.005 54.630 144.035 ;
        RECT 54.045 143.645 54.215 144.005 ;
        RECT 50.450 143.615 51.100 143.645 ;
        RECT 53.630 143.615 54.630 143.645 ;
        RECT 49.565 143.550 51.120 143.615 ;
        RECT 49.560 143.445 51.120 143.550 ;
        RECT 53.610 143.445 54.650 143.615 ;
        RECT 49.560 143.190 49.860 143.445 ;
        RECT 50.450 143.415 51.100 143.445 ;
        RECT 53.630 143.415 54.630 143.445 ;
        RECT 49.565 142.115 49.855 143.190 ;
        RECT 50.060 143.160 50.290 143.305 ;
        RECT 51.260 143.160 51.490 143.305 ;
        RECT 53.195 143.235 53.425 143.305 ;
        RECT 53.195 143.160 53.810 143.235 ;
        RECT 54.835 143.160 55.065 143.305 ;
        RECT 50.060 142.990 55.065 143.160 ;
        RECT 50.060 142.845 50.290 142.990 ;
        RECT 51.260 142.845 51.490 142.990 ;
        RECT 53.195 142.915 53.810 142.990 ;
        RECT 53.195 142.845 53.425 142.915 ;
        RECT 54.835 142.845 55.065 142.990 ;
        RECT 50.450 142.705 51.100 142.735 ;
        RECT 52.235 142.705 52.495 142.780 ;
        RECT 53.630 142.705 54.630 142.735 ;
        RECT 50.430 142.535 52.495 142.705 ;
        RECT 53.610 142.535 54.650 142.705 ;
        RECT 50.450 142.505 51.100 142.535 ;
        RECT 52.235 142.460 52.495 142.535 ;
        RECT 53.630 142.505 54.630 142.535 ;
        RECT 54.045 142.145 54.215 142.505 ;
        RECT 50.450 142.115 51.100 142.145 ;
        RECT 53.630 142.115 54.630 142.145 ;
        RECT 36.640 141.490 41.645 141.660 ;
        RECT 36.640 141.345 36.870 141.490 ;
        RECT 37.840 141.345 38.070 141.490 ;
        RECT 39.775 141.345 40.005 141.490 ;
        RECT 40.970 141.415 41.230 141.490 ;
        RECT 41.415 141.345 41.645 141.490 ;
        RECT 37.030 141.205 37.680 141.235 ;
        RECT 38.815 141.205 39.075 141.280 ;
        RECT 40.210 141.205 41.210 141.235 ;
        RECT 37.010 141.035 41.230 141.205 ;
        RECT 37.030 141.005 37.680 141.035 ;
        RECT 38.815 140.960 39.075 141.035 ;
        RECT 40.210 141.005 41.210 141.035 ;
        RECT 41.805 140.825 42.095 141.690 ;
        RECT 42.855 140.825 43.145 141.945 ;
        RECT 43.740 141.915 44.390 141.945 ;
        RECT 46.920 141.915 47.920 141.945 ;
        RECT 43.350 141.660 43.580 141.805 ;
        RECT 44.550 141.660 44.780 141.805 ;
        RECT 46.485 141.660 46.715 141.805 ;
        RECT 47.680 141.660 47.940 141.735 ;
        RECT 48.125 141.660 48.355 141.805 ;
        RECT 48.510 141.690 48.810 142.050 ;
        RECT 49.565 141.945 51.120 142.115 ;
        RECT 53.610 141.945 54.650 142.115 ;
        RECT 55.225 142.050 55.515 144.690 ;
        RECT 56.275 143.615 56.565 144.945 ;
        RECT 57.160 144.915 57.810 144.945 ;
        RECT 60.340 144.915 61.340 144.945 ;
        RECT 56.770 144.660 57.000 144.805 ;
        RECT 57.970 144.660 58.200 144.805 ;
        RECT 59.905 144.735 60.135 144.805 ;
        RECT 59.840 144.660 60.135 144.735 ;
        RECT 61.545 144.660 61.775 144.805 ;
        RECT 61.930 144.690 62.230 144.945 ;
        RECT 62.985 144.945 64.540 145.115 ;
        RECT 67.030 145.050 68.935 145.115 ;
        RECT 69.695 145.115 69.985 146.190 ;
        RECT 70.190 146.160 70.420 146.305 ;
        RECT 71.390 146.160 71.620 146.305 ;
        RECT 73.325 146.160 73.555 146.305 ;
        RECT 74.520 146.160 74.780 146.235 ;
        RECT 74.965 146.160 75.195 146.305 ;
        RECT 70.190 145.990 75.195 146.160 ;
        RECT 70.190 145.845 70.420 145.990 ;
        RECT 71.390 145.845 71.620 145.990 ;
        RECT 73.325 145.845 73.555 145.990 ;
        RECT 74.520 145.915 74.780 145.990 ;
        RECT 74.965 145.845 75.195 145.990 ;
        RECT 70.580 145.705 71.230 145.735 ;
        RECT 72.365 145.705 72.625 145.780 ;
        RECT 73.760 145.705 74.760 145.735 ;
        RECT 70.560 145.535 74.780 145.705 ;
        RECT 70.580 145.505 71.230 145.535 ;
        RECT 72.365 145.460 72.625 145.535 ;
        RECT 73.760 145.505 74.760 145.535 ;
        RECT 70.580 145.115 71.230 145.145 ;
        RECT 73.760 145.115 74.760 145.145 ;
        RECT 75.355 145.115 75.645 147.690 ;
        RECT 76.405 146.615 76.695 147.945 ;
        RECT 77.290 147.915 77.940 147.945 ;
        RECT 80.470 147.915 81.470 147.945 ;
        RECT 76.900 147.660 77.130 147.805 ;
        RECT 78.100 147.660 78.330 147.805 ;
        RECT 80.035 147.660 80.265 147.805 ;
        RECT 80.810 147.660 81.070 147.735 ;
        RECT 81.675 147.660 81.905 147.805 ;
        RECT 82.060 147.690 82.360 148.050 ;
        RECT 83.115 147.945 84.670 148.115 ;
        RECT 87.160 147.945 88.200 148.115 ;
        RECT 88.775 148.050 89.065 149.445 ;
        RECT 89.820 149.445 91.380 149.550 ;
        RECT 93.870 149.445 95.775 149.615 ;
        RECT 96.535 149.615 96.825 150.945 ;
        RECT 97.420 150.915 98.070 150.945 ;
        RECT 100.600 150.915 101.600 150.945 ;
        RECT 97.030 150.660 97.260 150.805 ;
        RECT 98.230 150.660 98.460 150.805 ;
        RECT 99.205 150.660 99.465 150.735 ;
        RECT 100.165 150.660 100.395 150.805 ;
        RECT 101.805 150.660 102.035 150.805 ;
        RECT 102.190 150.690 102.490 150.945 ;
        RECT 97.030 150.490 102.035 150.660 ;
        RECT 97.030 150.345 97.260 150.490 ;
        RECT 98.230 150.345 98.460 150.490 ;
        RECT 99.205 150.415 99.465 150.490 ;
        RECT 100.165 150.345 100.395 150.490 ;
        RECT 101.805 150.345 102.035 150.490 ;
        RECT 97.400 150.235 97.660 150.280 ;
        RECT 97.400 150.205 98.070 150.235 ;
        RECT 100.600 150.205 101.600 150.235 ;
        RECT 97.400 150.035 101.620 150.205 ;
        RECT 97.400 150.005 98.070 150.035 ;
        RECT 100.600 150.005 101.600 150.035 ;
        RECT 97.400 149.960 97.660 150.005 ;
        RECT 97.420 149.615 98.070 149.645 ;
        RECT 100.600 149.615 101.600 149.645 ;
        RECT 102.195 149.615 102.485 150.690 ;
        RECT 96.535 149.550 98.090 149.615 ;
        RECT 89.820 149.190 90.120 149.445 ;
        RECT 90.710 149.415 91.360 149.445 ;
        RECT 93.890 149.415 94.890 149.445 ;
        RECT 89.825 148.115 90.115 149.190 ;
        RECT 90.320 149.160 90.550 149.305 ;
        RECT 91.520 149.160 91.750 149.305 ;
        RECT 93.455 149.235 93.685 149.305 ;
        RECT 93.390 149.160 93.685 149.235 ;
        RECT 95.095 149.160 95.325 149.305 ;
        RECT 90.320 148.990 95.325 149.160 ;
        RECT 90.320 148.845 90.550 148.990 ;
        RECT 91.520 148.845 91.750 148.990 ;
        RECT 93.390 148.915 93.685 148.990 ;
        RECT 93.455 148.845 93.685 148.915 ;
        RECT 95.095 148.845 95.325 148.990 ;
        RECT 90.710 148.705 91.360 148.735 ;
        RECT 92.495 148.705 92.755 148.780 ;
        RECT 93.890 148.705 94.890 148.735 ;
        RECT 90.690 148.535 92.755 148.705 ;
        RECT 93.870 148.535 94.910 148.705 ;
        RECT 90.710 148.505 91.360 148.535 ;
        RECT 92.495 148.460 92.755 148.535 ;
        RECT 93.890 148.505 94.890 148.535 ;
        RECT 94.305 148.145 94.475 148.505 ;
        RECT 90.710 148.115 91.360 148.145 ;
        RECT 93.890 148.115 94.890 148.145 ;
        RECT 76.900 147.490 81.905 147.660 ;
        RECT 76.900 147.345 77.130 147.490 ;
        RECT 78.100 147.345 78.330 147.490 ;
        RECT 80.035 147.345 80.265 147.490 ;
        RECT 80.810 147.415 81.070 147.490 ;
        RECT 81.675 147.345 81.905 147.490 ;
        RECT 77.290 147.205 77.940 147.235 ;
        RECT 79.075 147.205 79.335 147.280 ;
        RECT 80.470 147.205 81.470 147.235 ;
        RECT 77.270 147.035 79.335 147.205 ;
        RECT 80.450 147.035 81.490 147.205 ;
        RECT 77.290 147.005 77.940 147.035 ;
        RECT 79.075 146.960 79.335 147.035 ;
        RECT 80.470 147.005 81.470 147.035 ;
        RECT 80.885 146.645 81.055 147.005 ;
        RECT 77.290 146.615 77.940 146.645 ;
        RECT 80.470 146.615 81.470 146.645 ;
        RECT 76.405 146.550 77.960 146.615 ;
        RECT 76.400 146.445 77.960 146.550 ;
        RECT 80.450 146.445 81.490 146.615 ;
        RECT 76.400 146.190 76.700 146.445 ;
        RECT 77.290 146.415 77.940 146.445 ;
        RECT 80.470 146.415 81.470 146.445 ;
        RECT 67.030 144.945 68.940 145.050 ;
        RECT 56.770 144.490 61.775 144.660 ;
        RECT 56.770 144.345 57.000 144.490 ;
        RECT 57.970 144.345 58.200 144.490 ;
        RECT 59.840 144.415 60.135 144.490 ;
        RECT 59.905 144.345 60.135 144.415 ;
        RECT 61.545 144.345 61.775 144.490 ;
        RECT 57.160 144.205 57.810 144.235 ;
        RECT 58.945 144.205 59.205 144.280 ;
        RECT 60.340 144.205 61.340 144.235 ;
        RECT 57.140 144.035 59.205 144.205 ;
        RECT 60.320 144.035 61.360 144.205 ;
        RECT 57.160 144.005 57.810 144.035 ;
        RECT 58.945 143.960 59.205 144.035 ;
        RECT 60.340 144.005 61.340 144.035 ;
        RECT 60.755 143.645 60.925 144.005 ;
        RECT 57.160 143.615 57.810 143.645 ;
        RECT 60.340 143.615 61.340 143.645 ;
        RECT 56.275 143.550 57.830 143.615 ;
        RECT 56.270 143.445 57.830 143.550 ;
        RECT 60.320 143.445 61.360 143.615 ;
        RECT 56.270 143.190 56.570 143.445 ;
        RECT 57.160 143.415 57.810 143.445 ;
        RECT 60.340 143.415 61.340 143.445 ;
        RECT 56.275 142.115 56.565 143.190 ;
        RECT 56.770 143.160 57.000 143.305 ;
        RECT 57.970 143.160 58.200 143.305 ;
        RECT 59.905 143.235 60.135 143.305 ;
        RECT 59.905 143.160 60.520 143.235 ;
        RECT 61.545 143.160 61.775 143.305 ;
        RECT 56.770 142.990 61.775 143.160 ;
        RECT 56.770 142.845 57.000 142.990 ;
        RECT 57.970 142.845 58.200 142.990 ;
        RECT 59.905 142.915 60.520 142.990 ;
        RECT 59.905 142.845 60.135 142.915 ;
        RECT 61.545 142.845 61.775 142.990 ;
        RECT 57.160 142.705 57.810 142.735 ;
        RECT 58.945 142.705 59.205 142.780 ;
        RECT 60.340 142.705 61.340 142.735 ;
        RECT 57.140 142.535 59.205 142.705 ;
        RECT 60.320 142.535 61.360 142.705 ;
        RECT 57.160 142.505 57.810 142.535 ;
        RECT 58.945 142.460 59.205 142.535 ;
        RECT 60.340 142.505 61.340 142.535 ;
        RECT 60.755 142.145 60.925 142.505 ;
        RECT 57.160 142.115 57.810 142.145 ;
        RECT 60.340 142.115 61.340 142.145 ;
        RECT 43.350 141.490 48.355 141.660 ;
        RECT 43.350 141.345 43.580 141.490 ;
        RECT 44.550 141.345 44.780 141.490 ;
        RECT 46.485 141.345 46.715 141.490 ;
        RECT 47.680 141.415 47.940 141.490 ;
        RECT 48.125 141.345 48.355 141.490 ;
        RECT 43.740 141.205 44.390 141.235 ;
        RECT 45.525 141.205 45.785 141.280 ;
        RECT 46.920 141.205 47.920 141.235 ;
        RECT 43.720 141.035 47.940 141.205 ;
        RECT 43.740 141.005 44.390 141.035 ;
        RECT 45.525 140.960 45.785 141.035 ;
        RECT 46.920 141.005 47.920 141.035 ;
        RECT 48.515 140.825 48.805 141.690 ;
        RECT 49.565 140.825 49.855 141.945 ;
        RECT 50.450 141.915 51.100 141.945 ;
        RECT 53.630 141.915 54.630 141.945 ;
        RECT 50.060 141.660 50.290 141.805 ;
        RECT 51.260 141.660 51.490 141.805 ;
        RECT 53.195 141.660 53.425 141.805 ;
        RECT 54.390 141.660 54.650 141.735 ;
        RECT 54.835 141.660 55.065 141.805 ;
        RECT 55.220 141.690 55.520 142.050 ;
        RECT 56.275 141.945 57.830 142.115 ;
        RECT 60.320 141.945 61.360 142.115 ;
        RECT 61.935 142.050 62.225 144.690 ;
        RECT 62.985 143.615 63.275 144.945 ;
        RECT 63.870 144.915 64.520 144.945 ;
        RECT 67.050 144.915 68.050 144.945 ;
        RECT 63.480 144.660 63.710 144.805 ;
        RECT 64.680 144.660 64.910 144.805 ;
        RECT 66.615 144.735 66.845 144.805 ;
        RECT 66.550 144.660 66.845 144.735 ;
        RECT 68.255 144.660 68.485 144.805 ;
        RECT 68.640 144.690 68.940 144.945 ;
        RECT 69.695 144.945 71.250 145.115 ;
        RECT 73.740 145.050 75.645 145.115 ;
        RECT 76.405 145.115 76.695 146.190 ;
        RECT 76.900 146.160 77.130 146.305 ;
        RECT 78.100 146.160 78.330 146.305 ;
        RECT 80.035 146.160 80.265 146.305 ;
        RECT 81.230 146.160 81.490 146.235 ;
        RECT 81.675 146.160 81.905 146.305 ;
        RECT 76.900 145.990 81.905 146.160 ;
        RECT 76.900 145.845 77.130 145.990 ;
        RECT 78.100 145.845 78.330 145.990 ;
        RECT 80.035 145.845 80.265 145.990 ;
        RECT 81.230 145.915 81.490 145.990 ;
        RECT 81.675 145.845 81.905 145.990 ;
        RECT 77.290 145.705 77.940 145.735 ;
        RECT 79.075 145.705 79.335 145.780 ;
        RECT 80.470 145.705 81.470 145.735 ;
        RECT 77.270 145.535 81.490 145.705 ;
        RECT 77.290 145.505 77.940 145.535 ;
        RECT 79.075 145.460 79.335 145.535 ;
        RECT 80.470 145.505 81.470 145.535 ;
        RECT 77.290 145.115 77.940 145.145 ;
        RECT 80.470 145.115 81.470 145.145 ;
        RECT 82.065 145.115 82.355 147.690 ;
        RECT 83.115 146.615 83.405 147.945 ;
        RECT 84.000 147.915 84.650 147.945 ;
        RECT 87.180 147.915 88.180 147.945 ;
        RECT 83.610 147.660 83.840 147.805 ;
        RECT 84.810 147.660 85.040 147.805 ;
        RECT 86.745 147.660 86.975 147.805 ;
        RECT 87.520 147.660 87.780 147.735 ;
        RECT 88.385 147.660 88.615 147.805 ;
        RECT 88.770 147.690 89.070 148.050 ;
        RECT 89.825 147.945 91.380 148.115 ;
        RECT 93.870 147.945 94.910 148.115 ;
        RECT 95.485 148.050 95.775 149.445 ;
        RECT 96.530 149.445 98.090 149.550 ;
        RECT 100.580 149.445 102.485 149.615 ;
        RECT 96.530 149.190 96.830 149.445 ;
        RECT 97.420 149.415 98.070 149.445 ;
        RECT 100.600 149.415 101.600 149.445 ;
        RECT 96.535 148.115 96.825 149.190 ;
        RECT 97.030 149.160 97.260 149.305 ;
        RECT 98.230 149.160 98.460 149.305 ;
        RECT 100.165 149.235 100.395 149.305 ;
        RECT 100.100 149.160 100.395 149.235 ;
        RECT 101.805 149.160 102.035 149.305 ;
        RECT 97.030 148.990 102.035 149.160 ;
        RECT 97.030 148.845 97.260 148.990 ;
        RECT 98.230 148.845 98.460 148.990 ;
        RECT 100.100 148.915 100.395 148.990 ;
        RECT 100.165 148.845 100.395 148.915 ;
        RECT 101.805 148.845 102.035 148.990 ;
        RECT 97.420 148.705 98.070 148.735 ;
        RECT 99.205 148.705 99.465 148.780 ;
        RECT 100.600 148.705 101.600 148.735 ;
        RECT 97.400 148.535 99.465 148.705 ;
        RECT 100.580 148.535 101.620 148.705 ;
        RECT 97.420 148.505 98.070 148.535 ;
        RECT 99.205 148.460 99.465 148.535 ;
        RECT 100.600 148.505 101.600 148.535 ;
        RECT 101.015 148.145 101.185 148.505 ;
        RECT 97.420 148.115 98.070 148.145 ;
        RECT 100.600 148.115 101.600 148.145 ;
        RECT 83.610 147.490 88.615 147.660 ;
        RECT 83.610 147.345 83.840 147.490 ;
        RECT 84.810 147.345 85.040 147.490 ;
        RECT 86.745 147.345 86.975 147.490 ;
        RECT 87.520 147.415 87.780 147.490 ;
        RECT 88.385 147.345 88.615 147.490 ;
        RECT 84.000 147.205 84.650 147.235 ;
        RECT 85.785 147.205 86.045 147.280 ;
        RECT 87.180 147.205 88.180 147.235 ;
        RECT 83.980 147.035 86.045 147.205 ;
        RECT 87.160 147.035 88.200 147.205 ;
        RECT 84.000 147.005 84.650 147.035 ;
        RECT 85.785 146.960 86.045 147.035 ;
        RECT 87.180 147.005 88.180 147.035 ;
        RECT 87.595 146.645 87.765 147.005 ;
        RECT 84.000 146.615 84.650 146.645 ;
        RECT 87.180 146.615 88.180 146.645 ;
        RECT 83.115 146.550 84.670 146.615 ;
        RECT 83.110 146.445 84.670 146.550 ;
        RECT 87.160 146.445 88.200 146.615 ;
        RECT 83.110 146.190 83.410 146.445 ;
        RECT 84.000 146.415 84.650 146.445 ;
        RECT 87.180 146.415 88.180 146.445 ;
        RECT 73.740 144.945 75.650 145.050 ;
        RECT 63.480 144.490 68.485 144.660 ;
        RECT 63.480 144.345 63.710 144.490 ;
        RECT 64.680 144.345 64.910 144.490 ;
        RECT 66.550 144.415 66.845 144.490 ;
        RECT 66.615 144.345 66.845 144.415 ;
        RECT 68.255 144.345 68.485 144.490 ;
        RECT 63.870 144.205 64.520 144.235 ;
        RECT 65.655 144.205 65.915 144.280 ;
        RECT 67.050 144.205 68.050 144.235 ;
        RECT 63.850 144.035 65.915 144.205 ;
        RECT 67.030 144.035 68.070 144.205 ;
        RECT 63.870 144.005 64.520 144.035 ;
        RECT 65.655 143.960 65.915 144.035 ;
        RECT 67.050 144.005 68.050 144.035 ;
        RECT 67.465 143.645 67.635 144.005 ;
        RECT 63.870 143.615 64.520 143.645 ;
        RECT 67.050 143.615 68.050 143.645 ;
        RECT 62.985 143.550 64.540 143.615 ;
        RECT 62.980 143.445 64.540 143.550 ;
        RECT 67.030 143.445 68.070 143.615 ;
        RECT 62.980 143.190 63.280 143.445 ;
        RECT 63.870 143.415 64.520 143.445 ;
        RECT 67.050 143.415 68.050 143.445 ;
        RECT 62.985 142.115 63.275 143.190 ;
        RECT 63.480 143.160 63.710 143.305 ;
        RECT 64.680 143.160 64.910 143.305 ;
        RECT 66.615 143.235 66.845 143.305 ;
        RECT 66.615 143.160 67.230 143.235 ;
        RECT 68.255 143.160 68.485 143.305 ;
        RECT 63.480 142.990 68.485 143.160 ;
        RECT 63.480 142.845 63.710 142.990 ;
        RECT 64.680 142.845 64.910 142.990 ;
        RECT 66.615 142.915 67.230 142.990 ;
        RECT 66.615 142.845 66.845 142.915 ;
        RECT 68.255 142.845 68.485 142.990 ;
        RECT 63.870 142.705 64.520 142.735 ;
        RECT 65.655 142.705 65.915 142.780 ;
        RECT 67.050 142.705 68.050 142.735 ;
        RECT 63.850 142.535 65.915 142.705 ;
        RECT 67.030 142.535 68.070 142.705 ;
        RECT 63.870 142.505 64.520 142.535 ;
        RECT 65.655 142.460 65.915 142.535 ;
        RECT 67.050 142.505 68.050 142.535 ;
        RECT 67.465 142.145 67.635 142.505 ;
        RECT 63.870 142.115 64.520 142.145 ;
        RECT 67.050 142.115 68.050 142.145 ;
        RECT 50.060 141.490 55.065 141.660 ;
        RECT 50.060 141.345 50.290 141.490 ;
        RECT 51.260 141.345 51.490 141.490 ;
        RECT 53.195 141.345 53.425 141.490 ;
        RECT 54.390 141.415 54.650 141.490 ;
        RECT 54.835 141.345 55.065 141.490 ;
        RECT 50.450 141.205 51.100 141.235 ;
        RECT 52.235 141.205 52.495 141.280 ;
        RECT 53.630 141.205 54.630 141.235 ;
        RECT 50.430 141.035 54.650 141.205 ;
        RECT 50.450 141.005 51.100 141.035 ;
        RECT 52.235 140.960 52.495 141.035 ;
        RECT 53.630 141.005 54.630 141.035 ;
        RECT 55.225 140.825 55.515 141.690 ;
        RECT 56.275 140.825 56.565 141.945 ;
        RECT 57.160 141.915 57.810 141.945 ;
        RECT 60.340 141.915 61.340 141.945 ;
        RECT 56.770 141.660 57.000 141.805 ;
        RECT 57.970 141.660 58.200 141.805 ;
        RECT 59.905 141.660 60.135 141.805 ;
        RECT 61.100 141.660 61.360 141.735 ;
        RECT 61.545 141.660 61.775 141.805 ;
        RECT 61.930 141.690 62.230 142.050 ;
        RECT 62.985 141.945 64.540 142.115 ;
        RECT 67.030 141.945 68.070 142.115 ;
        RECT 68.645 142.050 68.935 144.690 ;
        RECT 69.695 143.615 69.985 144.945 ;
        RECT 70.580 144.915 71.230 144.945 ;
        RECT 73.760 144.915 74.760 144.945 ;
        RECT 70.190 144.660 70.420 144.805 ;
        RECT 71.390 144.660 71.620 144.805 ;
        RECT 73.325 144.735 73.555 144.805 ;
        RECT 73.260 144.660 73.555 144.735 ;
        RECT 74.965 144.660 75.195 144.805 ;
        RECT 75.350 144.690 75.650 144.945 ;
        RECT 76.405 144.945 77.960 145.115 ;
        RECT 80.450 145.050 82.355 145.115 ;
        RECT 83.115 145.115 83.405 146.190 ;
        RECT 83.610 146.160 83.840 146.305 ;
        RECT 84.810 146.160 85.040 146.305 ;
        RECT 86.745 146.160 86.975 146.305 ;
        RECT 87.940 146.160 88.200 146.235 ;
        RECT 88.385 146.160 88.615 146.305 ;
        RECT 83.610 145.990 88.615 146.160 ;
        RECT 83.610 145.845 83.840 145.990 ;
        RECT 84.810 145.845 85.040 145.990 ;
        RECT 86.745 145.845 86.975 145.990 ;
        RECT 87.940 145.915 88.200 145.990 ;
        RECT 88.385 145.845 88.615 145.990 ;
        RECT 84.000 145.705 84.650 145.735 ;
        RECT 85.785 145.705 86.045 145.780 ;
        RECT 87.180 145.705 88.180 145.735 ;
        RECT 83.980 145.535 88.200 145.705 ;
        RECT 84.000 145.505 84.650 145.535 ;
        RECT 85.785 145.460 86.045 145.535 ;
        RECT 87.180 145.505 88.180 145.535 ;
        RECT 84.000 145.115 84.650 145.145 ;
        RECT 87.180 145.115 88.180 145.145 ;
        RECT 88.775 145.115 89.065 147.690 ;
        RECT 89.825 146.615 90.115 147.945 ;
        RECT 90.710 147.915 91.360 147.945 ;
        RECT 93.890 147.915 94.890 147.945 ;
        RECT 90.320 147.660 90.550 147.805 ;
        RECT 91.520 147.660 91.750 147.805 ;
        RECT 93.455 147.660 93.685 147.805 ;
        RECT 94.230 147.660 94.490 147.735 ;
        RECT 95.095 147.660 95.325 147.805 ;
        RECT 95.480 147.690 95.780 148.050 ;
        RECT 96.535 147.945 98.090 148.115 ;
        RECT 100.580 147.945 101.620 148.115 ;
        RECT 102.195 148.050 102.485 149.445 ;
        RECT 90.320 147.490 95.325 147.660 ;
        RECT 90.320 147.345 90.550 147.490 ;
        RECT 91.520 147.345 91.750 147.490 ;
        RECT 93.455 147.345 93.685 147.490 ;
        RECT 94.230 147.415 94.490 147.490 ;
        RECT 95.095 147.345 95.325 147.490 ;
        RECT 90.710 147.205 91.360 147.235 ;
        RECT 92.495 147.205 92.755 147.280 ;
        RECT 93.890 147.205 94.890 147.235 ;
        RECT 90.690 147.035 92.755 147.205 ;
        RECT 93.870 147.035 94.910 147.205 ;
        RECT 90.710 147.005 91.360 147.035 ;
        RECT 92.495 146.960 92.755 147.035 ;
        RECT 93.890 147.005 94.890 147.035 ;
        RECT 94.305 146.645 94.475 147.005 ;
        RECT 90.710 146.615 91.360 146.645 ;
        RECT 93.890 146.615 94.890 146.645 ;
        RECT 89.825 146.550 91.380 146.615 ;
        RECT 89.820 146.445 91.380 146.550 ;
        RECT 93.870 146.445 94.910 146.615 ;
        RECT 89.820 146.190 90.120 146.445 ;
        RECT 90.710 146.415 91.360 146.445 ;
        RECT 93.890 146.415 94.890 146.445 ;
        RECT 80.450 144.945 82.360 145.050 ;
        RECT 70.190 144.490 75.195 144.660 ;
        RECT 70.190 144.345 70.420 144.490 ;
        RECT 71.390 144.345 71.620 144.490 ;
        RECT 73.260 144.415 73.555 144.490 ;
        RECT 73.325 144.345 73.555 144.415 ;
        RECT 74.965 144.345 75.195 144.490 ;
        RECT 70.580 144.205 71.230 144.235 ;
        RECT 72.365 144.205 72.625 144.280 ;
        RECT 73.760 144.205 74.760 144.235 ;
        RECT 70.560 144.035 72.625 144.205 ;
        RECT 73.740 144.035 74.780 144.205 ;
        RECT 70.580 144.005 71.230 144.035 ;
        RECT 72.365 143.960 72.625 144.035 ;
        RECT 73.760 144.005 74.760 144.035 ;
        RECT 74.175 143.645 74.345 144.005 ;
        RECT 70.580 143.615 71.230 143.645 ;
        RECT 73.760 143.615 74.760 143.645 ;
        RECT 69.695 143.550 71.250 143.615 ;
        RECT 69.690 143.445 71.250 143.550 ;
        RECT 73.740 143.445 74.780 143.615 ;
        RECT 69.690 143.190 69.990 143.445 ;
        RECT 70.580 143.415 71.230 143.445 ;
        RECT 73.760 143.415 74.760 143.445 ;
        RECT 69.695 142.115 69.985 143.190 ;
        RECT 70.190 143.160 70.420 143.305 ;
        RECT 71.390 143.160 71.620 143.305 ;
        RECT 73.325 143.235 73.555 143.305 ;
        RECT 73.325 143.160 73.940 143.235 ;
        RECT 74.965 143.160 75.195 143.305 ;
        RECT 70.190 142.990 75.195 143.160 ;
        RECT 70.190 142.845 70.420 142.990 ;
        RECT 71.390 142.845 71.620 142.990 ;
        RECT 73.325 142.915 73.940 142.990 ;
        RECT 73.325 142.845 73.555 142.915 ;
        RECT 74.965 142.845 75.195 142.990 ;
        RECT 70.580 142.705 71.230 142.735 ;
        RECT 72.365 142.705 72.625 142.780 ;
        RECT 73.760 142.705 74.760 142.735 ;
        RECT 70.560 142.535 72.625 142.705 ;
        RECT 73.740 142.535 74.780 142.705 ;
        RECT 70.580 142.505 71.230 142.535 ;
        RECT 72.365 142.460 72.625 142.535 ;
        RECT 73.760 142.505 74.760 142.535 ;
        RECT 74.175 142.145 74.345 142.505 ;
        RECT 70.580 142.115 71.230 142.145 ;
        RECT 73.760 142.115 74.760 142.145 ;
        RECT 56.770 141.490 61.775 141.660 ;
        RECT 56.770 141.345 57.000 141.490 ;
        RECT 57.970 141.345 58.200 141.490 ;
        RECT 59.905 141.345 60.135 141.490 ;
        RECT 61.100 141.415 61.360 141.490 ;
        RECT 61.545 141.345 61.775 141.490 ;
        RECT 57.160 141.205 57.810 141.235 ;
        RECT 58.945 141.205 59.205 141.280 ;
        RECT 60.340 141.205 61.340 141.235 ;
        RECT 57.140 141.035 61.360 141.205 ;
        RECT 57.160 141.005 57.810 141.035 ;
        RECT 58.945 140.960 59.205 141.035 ;
        RECT 60.340 141.005 61.340 141.035 ;
        RECT 61.935 140.825 62.225 141.690 ;
        RECT 62.985 140.825 63.275 141.945 ;
        RECT 63.870 141.915 64.520 141.945 ;
        RECT 67.050 141.915 68.050 141.945 ;
        RECT 63.480 141.660 63.710 141.805 ;
        RECT 64.680 141.660 64.910 141.805 ;
        RECT 66.615 141.660 66.845 141.805 ;
        RECT 67.810 141.660 68.070 141.735 ;
        RECT 68.255 141.660 68.485 141.805 ;
        RECT 68.640 141.690 68.940 142.050 ;
        RECT 69.695 141.945 71.250 142.115 ;
        RECT 73.740 141.945 74.780 142.115 ;
        RECT 75.355 142.050 75.645 144.690 ;
        RECT 76.405 143.615 76.695 144.945 ;
        RECT 77.290 144.915 77.940 144.945 ;
        RECT 80.470 144.915 81.470 144.945 ;
        RECT 76.900 144.660 77.130 144.805 ;
        RECT 78.100 144.660 78.330 144.805 ;
        RECT 80.035 144.735 80.265 144.805 ;
        RECT 79.970 144.660 80.265 144.735 ;
        RECT 81.675 144.660 81.905 144.805 ;
        RECT 82.060 144.690 82.360 144.945 ;
        RECT 83.115 144.945 84.670 145.115 ;
        RECT 87.160 145.050 89.065 145.115 ;
        RECT 89.825 145.115 90.115 146.190 ;
        RECT 90.320 146.160 90.550 146.305 ;
        RECT 91.520 146.160 91.750 146.305 ;
        RECT 93.455 146.160 93.685 146.305 ;
        RECT 94.650 146.160 94.910 146.235 ;
        RECT 95.095 146.160 95.325 146.305 ;
        RECT 90.320 145.990 95.325 146.160 ;
        RECT 90.320 145.845 90.550 145.990 ;
        RECT 91.520 145.845 91.750 145.990 ;
        RECT 93.455 145.845 93.685 145.990 ;
        RECT 94.650 145.915 94.910 145.990 ;
        RECT 95.095 145.845 95.325 145.990 ;
        RECT 90.710 145.705 91.360 145.735 ;
        RECT 92.495 145.705 92.755 145.780 ;
        RECT 93.890 145.705 94.890 145.735 ;
        RECT 90.690 145.535 94.910 145.705 ;
        RECT 90.710 145.505 91.360 145.535 ;
        RECT 92.495 145.460 92.755 145.535 ;
        RECT 93.890 145.505 94.890 145.535 ;
        RECT 90.710 145.115 91.360 145.145 ;
        RECT 93.890 145.115 94.890 145.145 ;
        RECT 95.485 145.115 95.775 147.690 ;
        RECT 96.535 146.615 96.825 147.945 ;
        RECT 97.420 147.915 98.070 147.945 ;
        RECT 100.600 147.915 101.600 147.945 ;
        RECT 97.030 147.660 97.260 147.805 ;
        RECT 98.230 147.660 98.460 147.805 ;
        RECT 100.165 147.660 100.395 147.805 ;
        RECT 100.940 147.660 101.200 147.735 ;
        RECT 101.805 147.660 102.035 147.805 ;
        RECT 102.190 147.690 102.490 148.050 ;
        RECT 97.030 147.490 102.035 147.660 ;
        RECT 97.030 147.345 97.260 147.490 ;
        RECT 98.230 147.345 98.460 147.490 ;
        RECT 100.165 147.345 100.395 147.490 ;
        RECT 100.940 147.415 101.200 147.490 ;
        RECT 101.805 147.345 102.035 147.490 ;
        RECT 97.420 147.205 98.070 147.235 ;
        RECT 99.205 147.205 99.465 147.280 ;
        RECT 100.600 147.205 101.600 147.235 ;
        RECT 97.400 147.035 99.465 147.205 ;
        RECT 100.580 147.035 101.620 147.205 ;
        RECT 97.420 147.005 98.070 147.035 ;
        RECT 99.205 146.960 99.465 147.035 ;
        RECT 100.600 147.005 101.600 147.035 ;
        RECT 101.015 146.645 101.185 147.005 ;
        RECT 97.420 146.615 98.070 146.645 ;
        RECT 100.600 146.615 101.600 146.645 ;
        RECT 96.535 146.550 98.090 146.615 ;
        RECT 96.530 146.445 98.090 146.550 ;
        RECT 100.580 146.445 101.620 146.615 ;
        RECT 96.530 146.190 96.830 146.445 ;
        RECT 97.420 146.415 98.070 146.445 ;
        RECT 100.600 146.415 101.600 146.445 ;
        RECT 87.160 144.945 89.070 145.050 ;
        RECT 76.900 144.490 81.905 144.660 ;
        RECT 76.900 144.345 77.130 144.490 ;
        RECT 78.100 144.345 78.330 144.490 ;
        RECT 79.970 144.415 80.265 144.490 ;
        RECT 80.035 144.345 80.265 144.415 ;
        RECT 81.675 144.345 81.905 144.490 ;
        RECT 77.290 144.205 77.940 144.235 ;
        RECT 79.075 144.205 79.335 144.280 ;
        RECT 80.470 144.205 81.470 144.235 ;
        RECT 77.270 144.035 79.335 144.205 ;
        RECT 80.450 144.035 81.490 144.205 ;
        RECT 77.290 144.005 77.940 144.035 ;
        RECT 79.075 143.960 79.335 144.035 ;
        RECT 80.470 144.005 81.470 144.035 ;
        RECT 80.885 143.645 81.055 144.005 ;
        RECT 77.290 143.615 77.940 143.645 ;
        RECT 80.470 143.615 81.470 143.645 ;
        RECT 76.405 143.550 77.960 143.615 ;
        RECT 76.400 143.445 77.960 143.550 ;
        RECT 80.450 143.445 81.490 143.615 ;
        RECT 76.400 143.190 76.700 143.445 ;
        RECT 77.290 143.415 77.940 143.445 ;
        RECT 80.470 143.415 81.470 143.445 ;
        RECT 76.405 142.115 76.695 143.190 ;
        RECT 76.900 143.160 77.130 143.305 ;
        RECT 78.100 143.160 78.330 143.305 ;
        RECT 80.035 143.235 80.265 143.305 ;
        RECT 80.035 143.160 80.650 143.235 ;
        RECT 81.675 143.160 81.905 143.305 ;
        RECT 76.900 142.990 81.905 143.160 ;
        RECT 76.900 142.845 77.130 142.990 ;
        RECT 78.100 142.845 78.330 142.990 ;
        RECT 80.035 142.915 80.650 142.990 ;
        RECT 80.035 142.845 80.265 142.915 ;
        RECT 81.675 142.845 81.905 142.990 ;
        RECT 77.290 142.705 77.940 142.735 ;
        RECT 79.075 142.705 79.335 142.780 ;
        RECT 80.470 142.705 81.470 142.735 ;
        RECT 77.270 142.535 79.335 142.705 ;
        RECT 80.450 142.535 81.490 142.705 ;
        RECT 77.290 142.505 77.940 142.535 ;
        RECT 79.075 142.460 79.335 142.535 ;
        RECT 80.470 142.505 81.470 142.535 ;
        RECT 80.885 142.145 81.055 142.505 ;
        RECT 77.290 142.115 77.940 142.145 ;
        RECT 80.470 142.115 81.470 142.145 ;
        RECT 63.480 141.490 68.485 141.660 ;
        RECT 63.480 141.345 63.710 141.490 ;
        RECT 64.680 141.345 64.910 141.490 ;
        RECT 66.615 141.345 66.845 141.490 ;
        RECT 67.810 141.415 68.070 141.490 ;
        RECT 68.255 141.345 68.485 141.490 ;
        RECT 63.870 141.205 64.520 141.235 ;
        RECT 65.655 141.205 65.915 141.280 ;
        RECT 67.050 141.205 68.050 141.235 ;
        RECT 63.850 141.035 68.070 141.205 ;
        RECT 63.870 141.005 64.520 141.035 ;
        RECT 65.655 140.960 65.915 141.035 ;
        RECT 67.050 141.005 68.050 141.035 ;
        RECT 68.645 140.825 68.935 141.690 ;
        RECT 69.695 140.825 69.985 141.945 ;
        RECT 70.580 141.915 71.230 141.945 ;
        RECT 73.760 141.915 74.760 141.945 ;
        RECT 70.190 141.660 70.420 141.805 ;
        RECT 71.390 141.660 71.620 141.805 ;
        RECT 73.325 141.660 73.555 141.805 ;
        RECT 74.520 141.660 74.780 141.735 ;
        RECT 74.965 141.660 75.195 141.805 ;
        RECT 75.350 141.690 75.650 142.050 ;
        RECT 76.405 141.945 77.960 142.115 ;
        RECT 80.450 141.945 81.490 142.115 ;
        RECT 82.065 142.050 82.355 144.690 ;
        RECT 83.115 143.615 83.405 144.945 ;
        RECT 84.000 144.915 84.650 144.945 ;
        RECT 87.180 144.915 88.180 144.945 ;
        RECT 83.610 144.660 83.840 144.805 ;
        RECT 84.810 144.660 85.040 144.805 ;
        RECT 86.745 144.735 86.975 144.805 ;
        RECT 86.680 144.660 86.975 144.735 ;
        RECT 88.385 144.660 88.615 144.805 ;
        RECT 88.770 144.690 89.070 144.945 ;
        RECT 89.825 144.945 91.380 145.115 ;
        RECT 93.870 145.050 95.775 145.115 ;
        RECT 96.535 145.115 96.825 146.190 ;
        RECT 97.030 146.160 97.260 146.305 ;
        RECT 98.230 146.160 98.460 146.305 ;
        RECT 100.165 146.160 100.395 146.305 ;
        RECT 101.360 146.160 101.620 146.235 ;
        RECT 101.805 146.160 102.035 146.305 ;
        RECT 97.030 145.990 102.035 146.160 ;
        RECT 97.030 145.845 97.260 145.990 ;
        RECT 98.230 145.845 98.460 145.990 ;
        RECT 100.165 145.845 100.395 145.990 ;
        RECT 101.360 145.915 101.620 145.990 ;
        RECT 101.805 145.845 102.035 145.990 ;
        RECT 97.420 145.705 98.070 145.735 ;
        RECT 99.205 145.705 99.465 145.780 ;
        RECT 100.600 145.705 101.600 145.735 ;
        RECT 97.400 145.535 101.620 145.705 ;
        RECT 97.420 145.505 98.070 145.535 ;
        RECT 99.205 145.460 99.465 145.535 ;
        RECT 100.600 145.505 101.600 145.535 ;
        RECT 97.420 145.115 98.070 145.145 ;
        RECT 100.600 145.115 101.600 145.145 ;
        RECT 102.195 145.115 102.485 147.690 ;
        RECT 93.870 144.945 95.780 145.050 ;
        RECT 83.610 144.490 88.615 144.660 ;
        RECT 83.610 144.345 83.840 144.490 ;
        RECT 84.810 144.345 85.040 144.490 ;
        RECT 86.680 144.415 86.975 144.490 ;
        RECT 86.745 144.345 86.975 144.415 ;
        RECT 88.385 144.345 88.615 144.490 ;
        RECT 84.000 144.205 84.650 144.235 ;
        RECT 85.785 144.205 86.045 144.280 ;
        RECT 87.180 144.205 88.180 144.235 ;
        RECT 83.980 144.035 86.045 144.205 ;
        RECT 87.160 144.035 88.200 144.205 ;
        RECT 84.000 144.005 84.650 144.035 ;
        RECT 85.785 143.960 86.045 144.035 ;
        RECT 87.180 144.005 88.180 144.035 ;
        RECT 87.595 143.645 87.765 144.005 ;
        RECT 84.000 143.615 84.650 143.645 ;
        RECT 87.180 143.615 88.180 143.645 ;
        RECT 83.115 143.550 84.670 143.615 ;
        RECT 83.110 143.445 84.670 143.550 ;
        RECT 87.160 143.445 88.200 143.615 ;
        RECT 83.110 143.190 83.410 143.445 ;
        RECT 84.000 143.415 84.650 143.445 ;
        RECT 87.180 143.415 88.180 143.445 ;
        RECT 83.115 142.115 83.405 143.190 ;
        RECT 83.610 143.160 83.840 143.305 ;
        RECT 84.810 143.160 85.040 143.305 ;
        RECT 86.745 143.235 86.975 143.305 ;
        RECT 86.745 143.160 87.360 143.235 ;
        RECT 88.385 143.160 88.615 143.305 ;
        RECT 83.610 142.990 88.615 143.160 ;
        RECT 83.610 142.845 83.840 142.990 ;
        RECT 84.810 142.845 85.040 142.990 ;
        RECT 86.745 142.915 87.360 142.990 ;
        RECT 86.745 142.845 86.975 142.915 ;
        RECT 88.385 142.845 88.615 142.990 ;
        RECT 84.000 142.705 84.650 142.735 ;
        RECT 85.785 142.705 86.045 142.780 ;
        RECT 87.180 142.705 88.180 142.735 ;
        RECT 83.980 142.535 86.045 142.705 ;
        RECT 87.160 142.535 88.200 142.705 ;
        RECT 84.000 142.505 84.650 142.535 ;
        RECT 85.785 142.460 86.045 142.535 ;
        RECT 87.180 142.505 88.180 142.535 ;
        RECT 87.595 142.145 87.765 142.505 ;
        RECT 84.000 142.115 84.650 142.145 ;
        RECT 87.180 142.115 88.180 142.145 ;
        RECT 70.190 141.490 75.195 141.660 ;
        RECT 70.190 141.345 70.420 141.490 ;
        RECT 71.390 141.345 71.620 141.490 ;
        RECT 73.325 141.345 73.555 141.490 ;
        RECT 74.520 141.415 74.780 141.490 ;
        RECT 74.965 141.345 75.195 141.490 ;
        RECT 70.580 141.205 71.230 141.235 ;
        RECT 72.365 141.205 72.625 141.280 ;
        RECT 73.760 141.205 74.760 141.235 ;
        RECT 70.560 141.035 74.780 141.205 ;
        RECT 70.580 141.005 71.230 141.035 ;
        RECT 72.365 140.960 72.625 141.035 ;
        RECT 73.760 141.005 74.760 141.035 ;
        RECT 75.355 140.825 75.645 141.690 ;
        RECT 76.405 140.825 76.695 141.945 ;
        RECT 77.290 141.915 77.940 141.945 ;
        RECT 80.470 141.915 81.470 141.945 ;
        RECT 76.900 141.660 77.130 141.805 ;
        RECT 78.100 141.660 78.330 141.805 ;
        RECT 80.035 141.660 80.265 141.805 ;
        RECT 81.230 141.660 81.490 141.735 ;
        RECT 81.675 141.660 81.905 141.805 ;
        RECT 82.060 141.690 82.360 142.050 ;
        RECT 83.115 141.945 84.670 142.115 ;
        RECT 87.160 141.945 88.200 142.115 ;
        RECT 88.775 142.050 89.065 144.690 ;
        RECT 89.825 143.615 90.115 144.945 ;
        RECT 90.710 144.915 91.360 144.945 ;
        RECT 93.890 144.915 94.890 144.945 ;
        RECT 90.320 144.660 90.550 144.805 ;
        RECT 91.520 144.660 91.750 144.805 ;
        RECT 93.455 144.735 93.685 144.805 ;
        RECT 93.390 144.660 93.685 144.735 ;
        RECT 95.095 144.660 95.325 144.805 ;
        RECT 95.480 144.690 95.780 144.945 ;
        RECT 96.535 144.945 98.090 145.115 ;
        RECT 100.580 145.050 102.485 145.115 ;
        RECT 100.580 144.945 102.490 145.050 ;
        RECT 90.320 144.490 95.325 144.660 ;
        RECT 90.320 144.345 90.550 144.490 ;
        RECT 91.520 144.345 91.750 144.490 ;
        RECT 93.390 144.415 93.685 144.490 ;
        RECT 93.455 144.345 93.685 144.415 ;
        RECT 95.095 144.345 95.325 144.490 ;
        RECT 90.710 144.205 91.360 144.235 ;
        RECT 92.495 144.205 92.755 144.280 ;
        RECT 93.890 144.205 94.890 144.235 ;
        RECT 90.690 144.035 92.755 144.205 ;
        RECT 93.870 144.035 94.910 144.205 ;
        RECT 90.710 144.005 91.360 144.035 ;
        RECT 92.495 143.960 92.755 144.035 ;
        RECT 93.890 144.005 94.890 144.035 ;
        RECT 94.305 143.645 94.475 144.005 ;
        RECT 90.710 143.615 91.360 143.645 ;
        RECT 93.890 143.615 94.890 143.645 ;
        RECT 89.825 143.550 91.380 143.615 ;
        RECT 89.820 143.445 91.380 143.550 ;
        RECT 93.870 143.445 94.910 143.615 ;
        RECT 89.820 143.190 90.120 143.445 ;
        RECT 90.710 143.415 91.360 143.445 ;
        RECT 93.890 143.415 94.890 143.445 ;
        RECT 89.825 142.115 90.115 143.190 ;
        RECT 90.320 143.160 90.550 143.305 ;
        RECT 91.520 143.160 91.750 143.305 ;
        RECT 93.455 143.235 93.685 143.305 ;
        RECT 93.455 143.160 94.070 143.235 ;
        RECT 95.095 143.160 95.325 143.305 ;
        RECT 90.320 142.990 95.325 143.160 ;
        RECT 90.320 142.845 90.550 142.990 ;
        RECT 91.520 142.845 91.750 142.990 ;
        RECT 93.455 142.915 94.070 142.990 ;
        RECT 93.455 142.845 93.685 142.915 ;
        RECT 95.095 142.845 95.325 142.990 ;
        RECT 90.710 142.705 91.360 142.735 ;
        RECT 92.495 142.705 92.755 142.780 ;
        RECT 93.890 142.705 94.890 142.735 ;
        RECT 90.690 142.535 92.755 142.705 ;
        RECT 93.870 142.535 94.910 142.705 ;
        RECT 90.710 142.505 91.360 142.535 ;
        RECT 92.495 142.460 92.755 142.535 ;
        RECT 93.890 142.505 94.890 142.535 ;
        RECT 94.305 142.145 94.475 142.505 ;
        RECT 90.710 142.115 91.360 142.145 ;
        RECT 93.890 142.115 94.890 142.145 ;
        RECT 76.900 141.490 81.905 141.660 ;
        RECT 76.900 141.345 77.130 141.490 ;
        RECT 78.100 141.345 78.330 141.490 ;
        RECT 80.035 141.345 80.265 141.490 ;
        RECT 81.230 141.415 81.490 141.490 ;
        RECT 81.675 141.345 81.905 141.490 ;
        RECT 77.290 141.205 77.940 141.235 ;
        RECT 79.075 141.205 79.335 141.280 ;
        RECT 80.470 141.205 81.470 141.235 ;
        RECT 77.270 141.035 81.490 141.205 ;
        RECT 77.290 141.005 77.940 141.035 ;
        RECT 79.075 140.960 79.335 141.035 ;
        RECT 80.470 141.005 81.470 141.035 ;
        RECT 82.065 140.825 82.355 141.690 ;
        RECT 83.115 140.825 83.405 141.945 ;
        RECT 84.000 141.915 84.650 141.945 ;
        RECT 87.180 141.915 88.180 141.945 ;
        RECT 83.610 141.660 83.840 141.805 ;
        RECT 84.810 141.660 85.040 141.805 ;
        RECT 86.745 141.660 86.975 141.805 ;
        RECT 87.940 141.660 88.200 141.735 ;
        RECT 88.385 141.660 88.615 141.805 ;
        RECT 88.770 141.690 89.070 142.050 ;
        RECT 89.825 141.945 91.380 142.115 ;
        RECT 93.870 141.945 94.910 142.115 ;
        RECT 95.485 142.050 95.775 144.690 ;
        RECT 96.535 143.615 96.825 144.945 ;
        RECT 97.420 144.915 98.070 144.945 ;
        RECT 100.600 144.915 101.600 144.945 ;
        RECT 97.030 144.660 97.260 144.805 ;
        RECT 98.230 144.660 98.460 144.805 ;
        RECT 100.165 144.735 100.395 144.805 ;
        RECT 100.100 144.660 100.395 144.735 ;
        RECT 101.805 144.660 102.035 144.805 ;
        RECT 102.190 144.690 102.490 144.945 ;
        RECT 97.030 144.490 102.035 144.660 ;
        RECT 97.030 144.345 97.260 144.490 ;
        RECT 98.230 144.345 98.460 144.490 ;
        RECT 100.100 144.415 100.395 144.490 ;
        RECT 100.165 144.345 100.395 144.415 ;
        RECT 101.805 144.345 102.035 144.490 ;
        RECT 97.420 144.205 98.070 144.235 ;
        RECT 99.205 144.205 99.465 144.280 ;
        RECT 100.600 144.205 101.600 144.235 ;
        RECT 97.400 144.035 99.465 144.205 ;
        RECT 100.580 144.035 101.620 144.205 ;
        RECT 97.420 144.005 98.070 144.035 ;
        RECT 99.205 143.960 99.465 144.035 ;
        RECT 100.600 144.005 101.600 144.035 ;
        RECT 101.015 143.645 101.185 144.005 ;
        RECT 97.420 143.615 98.070 143.645 ;
        RECT 100.600 143.615 101.600 143.645 ;
        RECT 96.535 143.550 98.090 143.615 ;
        RECT 96.530 143.445 98.090 143.550 ;
        RECT 100.580 143.445 101.620 143.615 ;
        RECT 96.530 143.190 96.830 143.445 ;
        RECT 97.420 143.415 98.070 143.445 ;
        RECT 100.600 143.415 101.600 143.445 ;
        RECT 96.535 142.115 96.825 143.190 ;
        RECT 97.030 143.160 97.260 143.305 ;
        RECT 98.230 143.160 98.460 143.305 ;
        RECT 100.165 143.235 100.395 143.305 ;
        RECT 100.165 143.160 100.780 143.235 ;
        RECT 101.805 143.160 102.035 143.305 ;
        RECT 97.030 142.990 102.035 143.160 ;
        RECT 97.030 142.845 97.260 142.990 ;
        RECT 98.230 142.845 98.460 142.990 ;
        RECT 100.165 142.915 100.780 142.990 ;
        RECT 100.165 142.845 100.395 142.915 ;
        RECT 101.805 142.845 102.035 142.990 ;
        RECT 97.420 142.705 98.070 142.735 ;
        RECT 99.205 142.705 99.465 142.780 ;
        RECT 100.600 142.705 101.600 142.735 ;
        RECT 97.400 142.535 99.465 142.705 ;
        RECT 100.580 142.535 101.620 142.705 ;
        RECT 97.420 142.505 98.070 142.535 ;
        RECT 99.205 142.460 99.465 142.535 ;
        RECT 100.600 142.505 101.600 142.535 ;
        RECT 101.015 142.145 101.185 142.505 ;
        RECT 97.420 142.115 98.070 142.145 ;
        RECT 100.600 142.115 101.600 142.145 ;
        RECT 83.610 141.490 88.615 141.660 ;
        RECT 83.610 141.345 83.840 141.490 ;
        RECT 84.810 141.345 85.040 141.490 ;
        RECT 86.745 141.345 86.975 141.490 ;
        RECT 87.940 141.415 88.200 141.490 ;
        RECT 88.385 141.345 88.615 141.490 ;
        RECT 84.000 141.205 84.650 141.235 ;
        RECT 85.785 141.205 86.045 141.280 ;
        RECT 87.180 141.205 88.180 141.235 ;
        RECT 83.980 141.035 88.200 141.205 ;
        RECT 84.000 141.005 84.650 141.035 ;
        RECT 85.785 140.960 86.045 141.035 ;
        RECT 87.180 141.005 88.180 141.035 ;
        RECT 88.775 140.825 89.065 141.690 ;
        RECT 89.825 140.825 90.115 141.945 ;
        RECT 90.710 141.915 91.360 141.945 ;
        RECT 93.890 141.915 94.890 141.945 ;
        RECT 90.320 141.660 90.550 141.805 ;
        RECT 91.520 141.660 91.750 141.805 ;
        RECT 93.455 141.660 93.685 141.805 ;
        RECT 94.650 141.660 94.910 141.735 ;
        RECT 95.095 141.660 95.325 141.805 ;
        RECT 95.480 141.690 95.780 142.050 ;
        RECT 96.535 141.945 98.090 142.115 ;
        RECT 100.580 141.945 101.620 142.115 ;
        RECT 102.195 142.050 102.485 144.690 ;
        RECT 90.320 141.490 95.325 141.660 ;
        RECT 90.320 141.345 90.550 141.490 ;
        RECT 91.520 141.345 91.750 141.490 ;
        RECT 93.455 141.345 93.685 141.490 ;
        RECT 94.650 141.415 94.910 141.490 ;
        RECT 95.095 141.345 95.325 141.490 ;
        RECT 90.710 141.205 91.360 141.235 ;
        RECT 92.495 141.205 92.755 141.280 ;
        RECT 93.890 141.205 94.890 141.235 ;
        RECT 90.690 141.035 94.910 141.205 ;
        RECT 90.710 141.005 91.360 141.035 ;
        RECT 92.495 140.960 92.755 141.035 ;
        RECT 93.890 141.005 94.890 141.035 ;
        RECT 95.485 140.825 95.775 141.690 ;
        RECT 96.535 140.825 96.825 141.945 ;
        RECT 97.420 141.915 98.070 141.945 ;
        RECT 100.600 141.915 101.600 141.945 ;
        RECT 97.030 141.660 97.260 141.805 ;
        RECT 98.230 141.660 98.460 141.805 ;
        RECT 100.165 141.660 100.395 141.805 ;
        RECT 101.360 141.660 101.620 141.735 ;
        RECT 101.805 141.660 102.035 141.805 ;
        RECT 102.190 141.690 102.490 142.050 ;
        RECT 97.030 141.490 102.035 141.660 ;
        RECT 97.030 141.345 97.260 141.490 ;
        RECT 98.230 141.345 98.460 141.490 ;
        RECT 100.165 141.345 100.395 141.490 ;
        RECT 101.360 141.415 101.620 141.490 ;
        RECT 101.805 141.345 102.035 141.490 ;
        RECT 97.420 141.205 98.070 141.235 ;
        RECT 99.205 141.205 99.465 141.280 ;
        RECT 100.600 141.205 101.600 141.235 ;
        RECT 97.400 141.035 101.620 141.205 ;
        RECT 97.420 141.005 98.070 141.035 ;
        RECT 99.205 140.960 99.465 141.035 ;
        RECT 100.600 141.005 101.600 141.035 ;
        RECT 102.195 140.825 102.485 141.690 ;
        RECT 59.820 140.000 60.080 140.075 ;
        RECT 99.205 140.000 99.465 140.075 ;
        RECT 59.820 139.830 99.465 140.000 ;
        RECT 59.820 139.755 60.080 139.830 ;
        RECT 99.205 139.755 99.465 139.830 ;
        RECT 61.200 139.615 61.460 139.690 ;
        RECT 102.690 139.615 102.950 139.690 ;
        RECT 61.200 139.445 102.950 139.615 ;
        RECT 61.200 139.370 61.460 139.445 ;
        RECT 102.690 139.370 102.950 139.445 ;
        RECT 62.580 139.230 62.840 139.305 ;
        RECT 92.495 139.230 92.755 139.305 ;
        RECT 62.580 139.060 92.755 139.230 ;
        RECT 62.580 138.985 62.840 139.060 ;
        RECT 92.495 138.985 92.755 139.060 ;
        RECT 63.960 138.845 64.220 138.920 ;
        RECT 95.980 138.845 96.240 138.920 ;
        RECT 63.960 138.675 96.240 138.845 ;
        RECT 63.960 138.600 64.220 138.675 ;
        RECT 95.980 138.600 96.240 138.675 ;
        RECT 65.340 138.460 65.600 138.535 ;
        RECT 85.785 138.460 86.045 138.535 ;
        RECT 65.340 138.290 86.045 138.460 ;
        RECT 65.340 138.215 65.600 138.290 ;
        RECT 85.785 138.215 86.045 138.290 ;
        RECT 66.720 138.075 66.980 138.150 ;
        RECT 89.270 138.075 89.530 138.150 ;
        RECT 66.720 137.905 89.530 138.075 ;
        RECT 66.720 137.830 66.980 137.905 ;
        RECT 89.270 137.830 89.530 137.905 ;
        RECT 68.100 137.690 68.360 137.765 ;
        RECT 79.075 137.690 79.335 137.765 ;
        RECT 68.100 137.520 79.335 137.690 ;
        RECT 68.100 137.445 68.360 137.520 ;
        RECT 79.075 137.445 79.335 137.520 ;
        RECT 69.480 137.305 69.740 137.380 ;
        RECT 82.560 137.305 82.820 137.380 ;
        RECT 69.480 137.135 82.820 137.305 ;
        RECT 69.480 137.060 69.740 137.135 ;
        RECT 82.560 137.060 82.820 137.135 ;
        RECT 70.860 136.920 71.120 136.995 ;
        RECT 72.735 136.920 72.995 136.995 ;
        RECT 70.860 136.750 72.995 136.920 ;
        RECT 70.860 136.675 71.120 136.750 ;
        RECT 72.735 136.675 72.995 136.750 ;
        RECT 72.240 136.535 72.500 136.610 ;
        RECT 75.850 136.535 76.110 136.610 ;
        RECT 72.240 136.365 76.110 136.535 ;
        RECT 72.240 136.290 72.500 136.365 ;
        RECT 75.850 136.290 76.110 136.365 ;
        RECT 66.025 136.150 66.285 136.225 ;
        RECT 73.620 136.150 73.880 136.225 ;
        RECT 66.025 135.980 73.880 136.150 ;
        RECT 66.025 135.905 66.285 135.980 ;
        RECT 73.620 135.905 73.880 135.980 ;
        RECT 68.770 135.765 69.030 135.840 ;
        RECT 75.000 135.765 75.260 135.840 ;
        RECT 68.770 135.595 75.260 135.765 ;
        RECT 68.770 135.520 69.030 135.595 ;
        RECT 75.000 135.520 75.260 135.595 ;
        RECT 52.235 135.380 52.495 135.455 ;
        RECT 58.945 135.380 59.205 135.455 ;
        RECT 76.380 135.380 76.640 135.455 ;
        RECT 52.235 135.210 57.875 135.380 ;
        RECT 52.235 135.135 52.495 135.210 ;
        RECT 55.720 134.995 55.980 135.070 ;
        RECT 55.720 134.825 57.490 134.995 ;
        RECT 55.720 134.750 55.980 134.825 ;
        RECT 57.320 134.225 57.490 134.825 ;
        RECT 57.705 134.610 57.875 135.210 ;
        RECT 58.945 135.210 76.640 135.380 ;
        RECT 58.945 135.135 59.205 135.210 ;
        RECT 76.380 135.135 76.640 135.210 ;
        RECT 62.060 134.995 62.320 135.070 ;
        RECT 77.760 134.995 78.020 135.070 ;
        RECT 62.060 134.825 78.020 134.995 ;
        RECT 62.060 134.750 62.320 134.825 ;
        RECT 77.760 134.750 78.020 134.825 ;
        RECT 79.140 134.610 79.400 134.685 ;
        RECT 57.705 134.440 79.400 134.610 ;
        RECT 79.140 134.365 79.400 134.440 ;
        RECT 80.520 134.225 80.780 134.300 ;
        RECT 57.320 134.055 80.780 134.225 ;
        RECT 80.520 133.980 80.780 134.055 ;
        RECT 56.245 132.685 82.465 132.975 ;
        RECT 54.800 129.355 56.050 132.435 ;
        RECT 56.705 132.250 57.165 132.480 ;
        RECT 56.335 131.440 56.655 132.090 ;
        RECT 56.820 131.280 57.050 132.250 ;
        RECT 57.305 132.090 57.535 132.685 ;
        RECT 58.085 132.250 58.545 132.480 ;
        RECT 57.215 131.440 57.535 132.090 ;
        RECT 57.715 131.440 58.035 132.090 ;
        RECT 58.200 131.280 58.430 132.250 ;
        RECT 58.685 132.090 58.915 132.685 ;
        RECT 59.465 132.250 59.925 132.480 ;
        RECT 58.595 131.440 58.915 132.090 ;
        RECT 59.095 131.440 59.415 132.090 ;
        RECT 59.580 131.280 59.810 132.250 ;
        RECT 60.065 132.090 60.295 132.685 ;
        RECT 60.845 132.250 61.305 132.480 ;
        RECT 59.975 131.440 60.295 132.090 ;
        RECT 60.475 131.440 60.795 132.090 ;
        RECT 60.960 131.280 61.190 132.250 ;
        RECT 61.445 132.090 61.675 132.685 ;
        RECT 62.225 132.250 62.685 132.480 ;
        RECT 61.355 131.440 61.675 132.090 ;
        RECT 61.855 131.440 62.175 132.090 ;
        RECT 62.340 131.280 62.570 132.250 ;
        RECT 62.825 132.090 63.055 132.685 ;
        RECT 63.605 132.250 64.065 132.480 ;
        RECT 62.735 131.440 63.055 132.090 ;
        RECT 63.235 131.440 63.555 132.090 ;
        RECT 63.720 131.280 63.950 132.250 ;
        RECT 64.205 132.090 64.435 132.685 ;
        RECT 64.985 132.250 65.445 132.480 ;
        RECT 64.115 131.440 64.435 132.090 ;
        RECT 64.615 131.440 64.935 132.090 ;
        RECT 65.100 131.280 65.330 132.250 ;
        RECT 65.585 132.090 65.815 132.685 ;
        RECT 66.365 132.250 66.825 132.480 ;
        RECT 65.495 131.440 65.815 132.090 ;
        RECT 65.995 131.440 66.315 132.090 ;
        RECT 66.480 131.280 66.710 132.250 ;
        RECT 66.965 132.090 67.195 132.685 ;
        RECT 67.745 132.250 68.205 132.480 ;
        RECT 66.875 131.440 67.195 132.090 ;
        RECT 67.375 131.440 67.695 132.090 ;
        RECT 67.860 131.280 68.090 132.250 ;
        RECT 68.345 132.090 68.575 132.685 ;
        RECT 69.125 132.250 69.585 132.480 ;
        RECT 68.255 131.440 68.575 132.090 ;
        RECT 68.755 131.440 69.075 132.090 ;
        RECT 69.240 131.280 69.470 132.250 ;
        RECT 69.725 132.090 69.955 132.685 ;
        RECT 70.505 132.250 70.965 132.480 ;
        RECT 69.635 131.440 69.955 132.090 ;
        RECT 70.135 131.440 70.455 132.090 ;
        RECT 70.620 131.280 70.850 132.250 ;
        RECT 71.105 132.090 71.335 132.685 ;
        RECT 71.885 132.250 72.345 132.480 ;
        RECT 71.015 131.440 71.335 132.090 ;
        RECT 71.515 131.440 71.835 132.090 ;
        RECT 72.000 131.280 72.230 132.250 ;
        RECT 72.485 132.090 72.715 132.685 ;
        RECT 73.265 132.250 73.725 132.480 ;
        RECT 72.395 131.440 72.715 132.090 ;
        RECT 72.895 131.440 73.215 132.090 ;
        RECT 73.380 131.280 73.610 132.250 ;
        RECT 73.865 132.090 74.095 132.685 ;
        RECT 74.645 132.250 75.105 132.480 ;
        RECT 73.775 131.440 74.095 132.090 ;
        RECT 74.275 131.440 74.595 132.090 ;
        RECT 74.760 131.280 74.990 132.250 ;
        RECT 75.245 132.090 75.475 132.685 ;
        RECT 76.025 132.250 76.485 132.480 ;
        RECT 75.155 131.440 75.475 132.090 ;
        RECT 75.655 131.440 75.975 132.090 ;
        RECT 76.140 131.280 76.370 132.250 ;
        RECT 76.625 132.090 76.855 132.685 ;
        RECT 77.405 132.250 77.865 132.480 ;
        RECT 76.535 131.440 76.855 132.090 ;
        RECT 77.035 131.440 77.355 132.090 ;
        RECT 77.520 131.280 77.750 132.250 ;
        RECT 78.005 132.090 78.235 132.685 ;
        RECT 78.785 132.250 79.245 132.480 ;
        RECT 77.915 131.440 78.235 132.090 ;
        RECT 78.415 131.440 78.735 132.090 ;
        RECT 78.900 131.280 79.130 132.250 ;
        RECT 79.385 132.090 79.615 132.685 ;
        RECT 80.165 132.250 80.625 132.480 ;
        RECT 79.295 131.440 79.615 132.090 ;
        RECT 79.795 131.440 80.115 132.090 ;
        RECT 80.280 131.280 80.510 132.250 ;
        RECT 80.765 132.090 80.995 132.685 ;
        RECT 81.545 132.250 82.005 132.480 ;
        RECT 80.675 131.440 80.995 132.090 ;
        RECT 81.175 131.440 81.495 132.090 ;
        RECT 81.660 131.280 81.890 132.250 ;
        RECT 82.145 132.090 82.375 132.685 ;
        RECT 82.055 131.440 82.375 132.090 ;
        RECT 56.705 131.050 57.165 131.280 ;
        RECT 58.085 131.050 58.545 131.280 ;
        RECT 59.465 131.050 59.925 131.280 ;
        RECT 60.845 131.050 61.305 131.280 ;
        RECT 62.225 131.050 62.685 131.280 ;
        RECT 63.605 131.050 64.065 131.280 ;
        RECT 64.985 131.050 65.445 131.280 ;
        RECT 66.365 131.050 66.825 131.280 ;
        RECT 67.745 131.050 68.205 131.280 ;
        RECT 69.125 131.050 69.585 131.280 ;
        RECT 70.505 131.050 70.965 131.280 ;
        RECT 71.885 131.050 72.345 131.280 ;
        RECT 73.265 131.050 73.725 131.280 ;
        RECT 74.645 131.050 75.105 131.280 ;
        RECT 76.025 131.050 76.485 131.280 ;
        RECT 77.405 131.050 77.865 131.280 ;
        RECT 78.785 131.050 79.245 131.280 ;
        RECT 80.165 131.050 80.625 131.280 ;
        RECT 81.545 131.050 82.005 131.280 ;
        RECT 56.820 130.740 57.165 131.050 ;
        RECT 58.200 130.740 58.545 131.050 ;
        RECT 59.580 130.740 59.925 131.050 ;
        RECT 60.960 130.740 61.305 131.050 ;
        RECT 62.340 130.740 62.685 131.050 ;
        RECT 63.720 130.740 64.065 131.050 ;
        RECT 65.100 130.740 65.445 131.050 ;
        RECT 66.480 130.740 66.825 131.050 ;
        RECT 67.860 130.740 68.205 131.050 ;
        RECT 69.240 130.740 69.585 131.050 ;
        RECT 70.620 130.740 70.965 131.050 ;
        RECT 72.000 130.740 72.345 131.050 ;
        RECT 73.380 130.740 73.725 131.050 ;
        RECT 74.760 130.740 75.105 131.050 ;
        RECT 76.140 130.740 76.485 131.050 ;
        RECT 77.520 130.740 77.865 131.050 ;
        RECT 78.900 130.740 79.245 131.050 ;
        RECT 80.280 130.740 80.625 131.050 ;
        RECT 81.660 130.740 82.005 131.050 ;
        RECT 56.705 130.510 57.165 130.740 ;
        RECT 58.085 130.510 58.545 130.740 ;
        RECT 59.465 130.510 59.925 130.740 ;
        RECT 60.845 130.510 61.305 130.740 ;
        RECT 62.225 130.510 62.685 130.740 ;
        RECT 63.605 130.510 64.065 130.740 ;
        RECT 64.985 130.510 65.445 130.740 ;
        RECT 66.365 130.510 66.825 130.740 ;
        RECT 67.745 130.510 68.205 130.740 ;
        RECT 69.125 130.510 69.585 130.740 ;
        RECT 70.505 130.510 70.965 130.740 ;
        RECT 71.885 130.510 72.345 130.740 ;
        RECT 73.265 130.510 73.725 130.740 ;
        RECT 74.645 130.510 75.105 130.740 ;
        RECT 76.025 130.510 76.485 130.740 ;
        RECT 77.405 130.510 77.865 130.740 ;
        RECT 78.785 130.510 79.245 130.740 ;
        RECT 80.165 130.510 80.625 130.740 ;
        RECT 81.545 130.510 82.005 130.740 ;
        RECT 56.335 129.700 56.655 130.350 ;
        RECT 55.550 123.190 56.050 127.515 ;
        RECT 56.335 127.170 56.565 129.700 ;
        RECT 56.820 129.555 57.050 130.510 ;
        RECT 57.215 129.700 57.535 130.350 ;
        RECT 56.705 129.295 57.165 129.555 ;
        RECT 56.705 127.330 57.165 127.650 ;
        RECT 56.335 126.170 56.655 127.170 ;
        RECT 56.335 126.165 56.565 126.170 ;
        RECT 56.820 125.965 57.050 127.330 ;
        RECT 57.305 127.170 57.535 129.700 ;
        RECT 57.215 126.170 57.535 127.170 ;
        RECT 57.305 125.985 57.535 126.170 ;
        RECT 57.715 129.700 58.035 130.350 ;
        RECT 57.715 127.170 57.945 129.700 ;
        RECT 58.200 129.555 58.430 130.510 ;
        RECT 58.595 129.700 58.915 130.350 ;
        RECT 58.085 129.295 58.545 129.555 ;
        RECT 58.085 127.330 58.545 127.650 ;
        RECT 57.715 126.170 58.035 127.170 ;
        RECT 57.715 126.165 57.945 126.170 ;
        RECT 56.335 125.735 57.165 125.965 ;
        RECT 56.335 124.990 56.565 125.735 ;
        RECT 57.305 125.665 57.565 125.985 ;
        RECT 58.200 125.965 58.430 127.330 ;
        RECT 58.685 127.170 58.915 129.700 ;
        RECT 58.595 126.170 58.915 127.170 ;
        RECT 58.685 125.985 58.915 126.170 ;
        RECT 59.095 129.700 59.415 130.350 ;
        RECT 59.095 127.170 59.325 129.700 ;
        RECT 59.580 129.555 59.810 130.510 ;
        RECT 59.975 129.700 60.295 130.350 ;
        RECT 59.465 129.295 59.925 129.555 ;
        RECT 59.465 127.330 59.925 127.650 ;
        RECT 59.095 126.170 59.415 127.170 ;
        RECT 59.095 126.165 59.325 126.170 ;
        RECT 57.715 125.735 58.545 125.965 ;
        RECT 56.705 125.180 57.165 125.440 ;
        RECT 56.335 123.990 56.655 124.990 ;
        RECT 56.335 123.985 56.565 123.990 ;
        RECT 56.820 123.785 57.050 125.180 ;
        RECT 57.715 124.990 57.945 125.735 ;
        RECT 58.685 125.665 58.945 125.985 ;
        RECT 59.580 125.965 59.810 127.330 ;
        RECT 60.065 127.170 60.295 129.700 ;
        RECT 59.975 126.170 60.295 127.170 ;
        RECT 60.065 125.985 60.295 126.170 ;
        RECT 60.475 129.700 60.795 130.350 ;
        RECT 60.475 127.170 60.705 129.700 ;
        RECT 60.960 129.555 61.190 130.510 ;
        RECT 61.355 129.700 61.675 130.350 ;
        RECT 60.845 129.295 61.305 129.555 ;
        RECT 60.845 127.330 61.305 127.650 ;
        RECT 60.475 126.170 60.795 127.170 ;
        RECT 60.475 126.165 60.705 126.170 ;
        RECT 59.095 125.735 59.925 125.965 ;
        RECT 58.085 125.180 58.545 125.440 ;
        RECT 57.215 123.990 57.535 124.990 ;
        RECT 56.705 123.555 57.165 123.785 ;
        RECT 57.305 123.395 57.535 123.990 ;
        RECT 57.715 123.990 58.035 124.990 ;
        RECT 57.715 123.985 57.945 123.990 ;
        RECT 58.200 123.785 58.430 125.180 ;
        RECT 59.095 124.990 59.325 125.735 ;
        RECT 60.065 125.665 60.325 125.985 ;
        RECT 60.960 125.965 61.190 127.330 ;
        RECT 61.445 127.170 61.675 129.700 ;
        RECT 61.355 126.170 61.675 127.170 ;
        RECT 61.445 125.985 61.675 126.170 ;
        RECT 61.855 129.700 62.175 130.350 ;
        RECT 61.855 127.170 62.085 129.700 ;
        RECT 62.340 129.555 62.570 130.510 ;
        RECT 62.735 129.700 63.055 130.350 ;
        RECT 62.225 129.295 62.685 129.555 ;
        RECT 62.225 127.330 62.685 127.650 ;
        RECT 61.855 126.170 62.175 127.170 ;
        RECT 61.855 126.165 62.085 126.170 ;
        RECT 60.475 125.735 61.305 125.965 ;
        RECT 59.465 125.180 59.925 125.440 ;
        RECT 58.595 123.990 58.915 124.990 ;
        RECT 58.085 123.555 58.545 123.785 ;
        RECT 58.685 123.395 58.915 123.990 ;
        RECT 59.095 123.990 59.415 124.990 ;
        RECT 59.095 123.985 59.325 123.990 ;
        RECT 59.580 123.785 59.810 125.180 ;
        RECT 60.475 124.990 60.705 125.735 ;
        RECT 61.445 125.665 61.705 125.985 ;
        RECT 62.340 125.965 62.570 127.330 ;
        RECT 62.825 127.170 63.055 129.700 ;
        RECT 62.735 126.170 63.055 127.170 ;
        RECT 62.825 125.985 63.055 126.170 ;
        RECT 63.235 129.700 63.555 130.350 ;
        RECT 63.235 127.170 63.465 129.700 ;
        RECT 63.720 129.555 63.950 130.510 ;
        RECT 64.115 129.700 64.435 130.350 ;
        RECT 63.605 129.295 64.065 129.555 ;
        RECT 63.605 127.330 64.065 127.650 ;
        RECT 63.235 126.170 63.555 127.170 ;
        RECT 63.235 126.165 63.465 126.170 ;
        RECT 61.855 125.735 62.685 125.965 ;
        RECT 60.845 125.180 61.305 125.440 ;
        RECT 59.975 123.990 60.295 124.990 ;
        RECT 59.465 123.555 59.925 123.785 ;
        RECT 60.065 123.395 60.295 123.990 ;
        RECT 60.475 123.990 60.795 124.990 ;
        RECT 60.475 123.985 60.705 123.990 ;
        RECT 60.960 123.785 61.190 125.180 ;
        RECT 61.855 124.990 62.085 125.735 ;
        RECT 62.825 125.665 63.085 125.985 ;
        RECT 63.720 125.965 63.950 127.330 ;
        RECT 64.205 127.170 64.435 129.700 ;
        RECT 64.115 126.170 64.435 127.170 ;
        RECT 64.205 125.985 64.435 126.170 ;
        RECT 64.615 129.700 64.935 130.350 ;
        RECT 64.615 127.170 64.845 129.700 ;
        RECT 65.100 129.555 65.330 130.510 ;
        RECT 65.495 129.700 65.815 130.350 ;
        RECT 64.985 129.295 65.445 129.555 ;
        RECT 64.985 127.330 65.445 127.650 ;
        RECT 64.615 126.170 64.935 127.170 ;
        RECT 64.615 126.165 64.845 126.170 ;
        RECT 63.235 125.735 64.065 125.965 ;
        RECT 62.225 125.180 62.685 125.440 ;
        RECT 61.355 123.990 61.675 124.990 ;
        RECT 60.845 123.555 61.305 123.785 ;
        RECT 61.445 123.395 61.675 123.990 ;
        RECT 61.855 123.990 62.175 124.990 ;
        RECT 61.855 123.985 62.085 123.990 ;
        RECT 62.340 123.785 62.570 125.180 ;
        RECT 63.235 124.990 63.465 125.735 ;
        RECT 64.205 125.665 64.465 125.985 ;
        RECT 65.100 125.965 65.330 127.330 ;
        RECT 65.585 127.170 65.815 129.700 ;
        RECT 65.495 126.170 65.815 127.170 ;
        RECT 65.585 125.985 65.815 126.170 ;
        RECT 65.995 129.700 66.315 130.350 ;
        RECT 65.995 127.170 66.225 129.700 ;
        RECT 66.480 129.555 66.710 130.510 ;
        RECT 66.875 129.700 67.195 130.350 ;
        RECT 66.365 129.295 66.825 129.555 ;
        RECT 66.365 127.330 66.825 127.650 ;
        RECT 65.995 126.170 66.315 127.170 ;
        RECT 65.995 126.165 66.225 126.170 ;
        RECT 64.615 125.735 65.445 125.965 ;
        RECT 63.605 125.180 64.065 125.440 ;
        RECT 62.735 123.990 63.055 124.990 ;
        RECT 62.225 123.555 62.685 123.785 ;
        RECT 62.825 123.395 63.055 123.990 ;
        RECT 63.235 123.990 63.555 124.990 ;
        RECT 63.235 123.985 63.465 123.990 ;
        RECT 63.720 123.785 63.950 125.180 ;
        RECT 64.615 124.990 64.845 125.735 ;
        RECT 65.585 125.665 65.845 125.985 ;
        RECT 66.480 125.965 66.710 127.330 ;
        RECT 66.965 127.170 67.195 129.700 ;
        RECT 66.875 126.170 67.195 127.170 ;
        RECT 66.965 125.985 67.195 126.170 ;
        RECT 67.375 129.700 67.695 130.350 ;
        RECT 67.375 127.170 67.605 129.700 ;
        RECT 67.860 129.555 68.090 130.510 ;
        RECT 68.255 129.700 68.575 130.350 ;
        RECT 67.745 129.295 68.205 129.555 ;
        RECT 67.745 127.330 68.205 127.650 ;
        RECT 67.375 126.170 67.695 127.170 ;
        RECT 67.375 126.165 67.605 126.170 ;
        RECT 65.995 125.735 66.825 125.965 ;
        RECT 64.985 125.180 65.445 125.440 ;
        RECT 64.115 123.990 64.435 124.990 ;
        RECT 63.605 123.555 64.065 123.785 ;
        RECT 64.205 123.395 64.435 123.990 ;
        RECT 64.615 123.990 64.935 124.990 ;
        RECT 64.615 123.985 64.845 123.990 ;
        RECT 65.100 123.785 65.330 125.180 ;
        RECT 65.995 124.990 66.225 125.735 ;
        RECT 66.965 125.665 67.225 125.985 ;
        RECT 67.860 125.965 68.090 127.330 ;
        RECT 68.345 127.170 68.575 129.700 ;
        RECT 68.255 126.170 68.575 127.170 ;
        RECT 68.345 125.985 68.575 126.170 ;
        RECT 68.755 129.700 69.075 130.350 ;
        RECT 68.755 127.170 68.985 129.700 ;
        RECT 69.240 129.555 69.470 130.510 ;
        RECT 69.635 129.700 69.955 130.350 ;
        RECT 69.125 129.295 69.585 129.555 ;
        RECT 69.125 127.330 69.585 127.650 ;
        RECT 68.755 126.170 69.075 127.170 ;
        RECT 68.755 126.165 68.985 126.170 ;
        RECT 67.375 125.735 68.205 125.965 ;
        RECT 66.365 125.180 66.825 125.440 ;
        RECT 65.495 123.990 65.815 124.990 ;
        RECT 64.985 123.555 65.445 123.785 ;
        RECT 65.585 123.395 65.815 123.990 ;
        RECT 65.995 123.990 66.315 124.990 ;
        RECT 65.995 123.985 66.225 123.990 ;
        RECT 66.480 123.785 66.710 125.180 ;
        RECT 67.375 124.990 67.605 125.735 ;
        RECT 68.345 125.665 68.605 125.985 ;
        RECT 69.240 125.965 69.470 127.330 ;
        RECT 69.725 127.170 69.955 129.700 ;
        RECT 69.635 126.170 69.955 127.170 ;
        RECT 69.725 125.985 69.955 126.170 ;
        RECT 70.135 129.700 70.455 130.350 ;
        RECT 70.135 127.170 70.365 129.700 ;
        RECT 70.620 129.555 70.850 130.510 ;
        RECT 71.015 129.700 71.335 130.350 ;
        RECT 70.505 129.295 70.965 129.555 ;
        RECT 70.505 127.330 70.965 127.650 ;
        RECT 70.135 126.170 70.455 127.170 ;
        RECT 70.135 126.165 70.365 126.170 ;
        RECT 68.755 125.735 69.585 125.965 ;
        RECT 67.745 125.180 68.205 125.440 ;
        RECT 66.875 123.990 67.195 124.990 ;
        RECT 66.365 123.555 66.825 123.785 ;
        RECT 66.965 123.395 67.195 123.990 ;
        RECT 67.375 123.990 67.695 124.990 ;
        RECT 67.375 123.985 67.605 123.990 ;
        RECT 67.860 123.785 68.090 125.180 ;
        RECT 68.755 124.990 68.985 125.735 ;
        RECT 69.725 125.665 69.985 125.985 ;
        RECT 70.620 125.965 70.850 127.330 ;
        RECT 71.105 127.170 71.335 129.700 ;
        RECT 71.015 126.170 71.335 127.170 ;
        RECT 71.105 125.985 71.335 126.170 ;
        RECT 71.515 129.700 71.835 130.350 ;
        RECT 71.515 127.170 71.745 129.700 ;
        RECT 72.000 129.555 72.230 130.510 ;
        RECT 72.395 129.700 72.715 130.350 ;
        RECT 71.885 129.295 72.345 129.555 ;
        RECT 71.885 127.330 72.345 127.650 ;
        RECT 71.515 126.170 71.835 127.170 ;
        RECT 71.515 126.165 71.745 126.170 ;
        RECT 70.135 125.735 70.965 125.965 ;
        RECT 69.125 125.180 69.585 125.440 ;
        RECT 68.255 123.990 68.575 124.990 ;
        RECT 67.745 123.555 68.205 123.785 ;
        RECT 68.345 123.395 68.575 123.990 ;
        RECT 68.755 123.990 69.075 124.990 ;
        RECT 68.755 123.985 68.985 123.990 ;
        RECT 69.240 123.785 69.470 125.180 ;
        RECT 70.135 124.990 70.365 125.735 ;
        RECT 71.105 125.665 71.365 125.985 ;
        RECT 72.000 125.965 72.230 127.330 ;
        RECT 72.485 127.170 72.715 129.700 ;
        RECT 72.395 126.170 72.715 127.170 ;
        RECT 72.485 125.985 72.715 126.170 ;
        RECT 72.895 129.700 73.215 130.350 ;
        RECT 72.895 127.170 73.125 129.700 ;
        RECT 73.380 129.555 73.610 130.510 ;
        RECT 73.775 129.700 74.095 130.350 ;
        RECT 73.265 129.295 73.725 129.555 ;
        RECT 73.265 127.330 73.725 127.650 ;
        RECT 72.895 126.170 73.215 127.170 ;
        RECT 72.895 126.165 73.125 126.170 ;
        RECT 71.515 125.735 72.345 125.965 ;
        RECT 70.505 125.180 70.965 125.440 ;
        RECT 69.635 123.990 69.955 124.990 ;
        RECT 69.125 123.555 69.585 123.785 ;
        RECT 69.725 123.395 69.955 123.990 ;
        RECT 70.135 123.990 70.455 124.990 ;
        RECT 70.135 123.985 70.365 123.990 ;
        RECT 70.620 123.785 70.850 125.180 ;
        RECT 71.515 124.990 71.745 125.735 ;
        RECT 72.485 125.665 72.745 125.985 ;
        RECT 73.380 125.965 73.610 127.330 ;
        RECT 73.865 127.170 74.095 129.700 ;
        RECT 73.775 126.170 74.095 127.170 ;
        RECT 73.865 125.985 74.095 126.170 ;
        RECT 74.275 129.700 74.595 130.350 ;
        RECT 74.275 127.170 74.505 129.700 ;
        RECT 74.760 129.555 74.990 130.510 ;
        RECT 75.155 129.700 75.475 130.350 ;
        RECT 74.645 129.295 75.105 129.555 ;
        RECT 74.645 127.330 75.105 127.650 ;
        RECT 74.275 126.170 74.595 127.170 ;
        RECT 74.275 126.165 74.505 126.170 ;
        RECT 72.895 125.735 73.725 125.965 ;
        RECT 71.885 125.180 72.345 125.440 ;
        RECT 71.015 123.990 71.335 124.990 ;
        RECT 70.505 123.555 70.965 123.785 ;
        RECT 71.105 123.395 71.335 123.990 ;
        RECT 71.515 123.990 71.835 124.990 ;
        RECT 71.515 123.985 71.745 123.990 ;
        RECT 72.000 123.785 72.230 125.180 ;
        RECT 72.895 124.990 73.125 125.735 ;
        RECT 73.865 125.665 74.125 125.985 ;
        RECT 74.760 125.965 74.990 127.330 ;
        RECT 75.245 127.170 75.475 129.700 ;
        RECT 75.155 126.170 75.475 127.170 ;
        RECT 75.245 125.985 75.475 126.170 ;
        RECT 75.655 129.700 75.975 130.350 ;
        RECT 75.655 127.170 75.885 129.700 ;
        RECT 76.140 129.555 76.370 130.510 ;
        RECT 76.535 129.700 76.855 130.350 ;
        RECT 76.025 129.295 76.485 129.555 ;
        RECT 76.025 127.330 76.485 127.650 ;
        RECT 75.655 126.170 75.975 127.170 ;
        RECT 75.655 126.165 75.885 126.170 ;
        RECT 74.275 125.735 75.105 125.965 ;
        RECT 73.265 125.180 73.725 125.440 ;
        RECT 72.395 123.990 72.715 124.990 ;
        RECT 71.885 123.555 72.345 123.785 ;
        RECT 72.485 123.395 72.715 123.990 ;
        RECT 72.895 123.990 73.215 124.990 ;
        RECT 72.895 123.985 73.125 123.990 ;
        RECT 73.380 123.785 73.610 125.180 ;
        RECT 74.275 124.990 74.505 125.735 ;
        RECT 75.245 125.665 75.505 125.985 ;
        RECT 76.140 125.965 76.370 127.330 ;
        RECT 76.625 127.170 76.855 129.700 ;
        RECT 76.535 126.170 76.855 127.170 ;
        RECT 76.625 125.985 76.855 126.170 ;
        RECT 77.035 129.700 77.355 130.350 ;
        RECT 77.035 127.170 77.265 129.700 ;
        RECT 77.520 129.555 77.750 130.510 ;
        RECT 77.915 129.700 78.235 130.350 ;
        RECT 77.405 129.295 77.865 129.555 ;
        RECT 77.405 127.330 77.865 127.650 ;
        RECT 77.035 126.170 77.355 127.170 ;
        RECT 77.035 126.165 77.265 126.170 ;
        RECT 75.655 125.735 76.485 125.965 ;
        RECT 74.645 125.180 75.105 125.440 ;
        RECT 73.775 123.990 74.095 124.990 ;
        RECT 73.265 123.555 73.725 123.785 ;
        RECT 73.865 123.395 74.095 123.990 ;
        RECT 74.275 123.990 74.595 124.990 ;
        RECT 74.275 123.985 74.505 123.990 ;
        RECT 74.760 123.785 74.990 125.180 ;
        RECT 75.655 124.990 75.885 125.735 ;
        RECT 76.625 125.665 76.885 125.985 ;
        RECT 77.520 125.965 77.750 127.330 ;
        RECT 78.005 127.170 78.235 129.700 ;
        RECT 77.915 126.170 78.235 127.170 ;
        RECT 78.005 125.985 78.235 126.170 ;
        RECT 78.415 129.700 78.735 130.350 ;
        RECT 78.415 127.170 78.645 129.700 ;
        RECT 78.900 129.555 79.130 130.510 ;
        RECT 79.295 129.700 79.615 130.350 ;
        RECT 78.785 129.295 79.245 129.555 ;
        RECT 78.785 127.330 79.245 127.650 ;
        RECT 78.415 126.170 78.735 127.170 ;
        RECT 78.415 126.165 78.645 126.170 ;
        RECT 77.035 125.735 77.865 125.965 ;
        RECT 76.025 125.180 76.485 125.440 ;
        RECT 75.155 123.990 75.475 124.990 ;
        RECT 74.645 123.555 75.105 123.785 ;
        RECT 75.245 123.395 75.475 123.990 ;
        RECT 75.655 123.990 75.975 124.990 ;
        RECT 75.655 123.985 75.885 123.990 ;
        RECT 76.140 123.785 76.370 125.180 ;
        RECT 77.035 124.990 77.265 125.735 ;
        RECT 78.005 125.665 78.265 125.985 ;
        RECT 78.900 125.965 79.130 127.330 ;
        RECT 79.385 127.170 79.615 129.700 ;
        RECT 79.295 126.170 79.615 127.170 ;
        RECT 79.385 125.985 79.615 126.170 ;
        RECT 79.795 129.700 80.115 130.350 ;
        RECT 79.795 127.170 80.025 129.700 ;
        RECT 80.280 129.555 80.510 130.510 ;
        RECT 80.675 129.700 80.995 130.350 ;
        RECT 80.165 129.295 80.625 129.555 ;
        RECT 80.165 127.330 80.625 127.650 ;
        RECT 79.795 126.170 80.115 127.170 ;
        RECT 79.795 126.165 80.025 126.170 ;
        RECT 78.415 125.735 79.245 125.965 ;
        RECT 77.405 125.180 77.865 125.440 ;
        RECT 76.535 123.990 76.855 124.990 ;
        RECT 76.025 123.555 76.485 123.785 ;
        RECT 76.625 123.395 76.855 123.990 ;
        RECT 77.035 123.990 77.355 124.990 ;
        RECT 77.035 123.985 77.265 123.990 ;
        RECT 77.520 123.785 77.750 125.180 ;
        RECT 78.415 124.990 78.645 125.735 ;
        RECT 79.385 125.665 79.645 125.985 ;
        RECT 80.280 125.965 80.510 127.330 ;
        RECT 80.765 127.170 80.995 129.700 ;
        RECT 80.675 126.170 80.995 127.170 ;
        RECT 80.765 125.985 80.995 126.170 ;
        RECT 81.175 129.700 81.495 130.350 ;
        RECT 81.175 127.170 81.405 129.700 ;
        RECT 81.660 129.555 81.890 130.510 ;
        RECT 82.055 129.700 82.375 130.350 ;
        RECT 81.545 129.295 82.005 129.555 ;
        RECT 81.545 127.330 82.005 127.650 ;
        RECT 81.175 126.170 81.495 127.170 ;
        RECT 81.175 126.165 81.405 126.170 ;
        RECT 79.795 125.735 80.625 125.965 ;
        RECT 78.785 125.180 79.245 125.440 ;
        RECT 77.915 123.990 78.235 124.990 ;
        RECT 77.405 123.555 77.865 123.785 ;
        RECT 78.005 123.395 78.235 123.990 ;
        RECT 78.415 123.990 78.735 124.990 ;
        RECT 78.415 123.985 78.645 123.990 ;
        RECT 78.900 123.785 79.130 125.180 ;
        RECT 79.795 124.990 80.025 125.735 ;
        RECT 80.765 125.665 81.025 125.985 ;
        RECT 81.660 125.965 81.890 127.330 ;
        RECT 82.145 127.170 82.375 129.700 ;
        RECT 82.660 129.355 83.910 132.435 ;
        RECT 82.055 126.170 82.375 127.170 ;
        RECT 82.145 125.985 82.375 126.170 ;
        RECT 81.175 125.735 82.005 125.965 ;
        RECT 80.165 125.180 80.625 125.440 ;
        RECT 79.295 123.990 79.615 124.990 ;
        RECT 78.785 123.555 79.245 123.785 ;
        RECT 79.385 123.395 79.615 123.990 ;
        RECT 79.795 123.990 80.115 124.990 ;
        RECT 79.795 123.985 80.025 123.990 ;
        RECT 80.280 123.785 80.510 125.180 ;
        RECT 81.175 124.990 81.405 125.735 ;
        RECT 82.145 125.665 82.405 125.985 ;
        RECT 81.545 125.180 82.005 125.440 ;
        RECT 80.675 123.990 80.995 124.990 ;
        RECT 80.165 123.555 80.625 123.785 ;
        RECT 80.765 123.395 80.995 123.990 ;
        RECT 81.175 123.990 81.495 124.990 ;
        RECT 81.175 123.985 81.405 123.990 ;
        RECT 81.660 123.785 81.890 125.180 ;
        RECT 82.055 123.990 82.375 124.990 ;
        RECT 81.545 123.555 82.005 123.785 ;
        RECT 82.145 123.395 82.375 123.990 ;
        RECT 56.245 123.105 82.465 123.395 ;
        RECT 82.660 123.190 83.160 127.515 ;
        RECT 54.800 121.120 55.360 121.350 ;
        RECT 83.350 121.120 83.910 121.350 ;
        RECT 54.800 118.960 57.080 121.120 ;
        RECT 57.560 118.960 58.740 121.120 ;
        RECT 59.220 118.960 60.400 121.120 ;
        RECT 60.880 118.960 62.060 121.120 ;
        RECT 62.540 118.960 63.720 121.120 ;
        RECT 64.200 118.960 65.380 121.120 ;
        RECT 65.860 118.960 67.040 121.120 ;
        RECT 67.520 118.960 68.700 121.120 ;
        RECT 54.800 110.370 55.360 118.960 ;
        RECT 69.180 113.540 69.530 121.120 ;
        RECT 70.010 118.360 70.360 121.120 ;
        RECT 70.840 118.960 72.020 121.120 ;
        RECT 72.500 118.960 73.680 121.120 ;
        RECT 74.160 118.960 75.340 121.120 ;
        RECT 75.820 118.960 77.000 121.120 ;
        RECT 77.480 118.960 78.660 121.120 ;
        RECT 79.140 118.960 80.320 121.120 ;
        RECT 80.800 118.960 81.980 121.120 ;
        RECT 82.460 118.960 83.910 121.120 ;
        RECT 69.150 113.190 69.560 113.540 ;
        RECT 83.350 110.370 83.910 118.960 ;
        RECT 54.800 108.210 56.250 110.370 ;
        RECT 56.730 108.210 57.910 110.370 ;
        RECT 58.390 108.210 59.570 110.370 ;
        RECT 60.050 108.210 61.230 110.370 ;
        RECT 61.710 108.210 62.890 110.370 ;
        RECT 63.370 108.210 64.550 110.370 ;
        RECT 65.030 108.210 66.210 110.370 ;
        RECT 66.690 108.210 67.870 110.370 ;
        RECT 68.350 108.210 69.530 110.370 ;
        RECT 70.010 108.210 71.190 110.370 ;
        RECT 71.670 108.210 72.850 110.370 ;
        RECT 73.330 108.210 74.510 110.370 ;
        RECT 74.990 108.210 76.170 110.370 ;
        RECT 76.650 108.210 77.830 110.370 ;
        RECT 78.310 108.210 79.490 110.370 ;
        RECT 79.970 108.210 81.150 110.370 ;
        RECT 81.630 108.210 81.980 110.370 ;
        RECT 82.460 108.210 83.910 110.370 ;
        RECT 54.800 107.980 55.360 108.210 ;
        RECT 83.350 107.980 83.910 108.210 ;
        RECT 55.550 101.815 56.050 106.140 ;
        RECT 56.245 105.935 82.465 106.225 ;
        RECT 56.335 105.340 56.565 105.935 ;
        RECT 56.705 105.545 57.165 105.775 ;
        RECT 56.335 104.340 56.655 105.340 ;
        RECT 56.820 104.150 57.050 105.545 ;
        RECT 57.305 105.340 57.535 105.345 ;
        RECT 57.215 104.340 57.535 105.340 ;
        RECT 57.715 105.340 57.945 105.935 ;
        RECT 58.085 105.545 58.545 105.775 ;
        RECT 57.715 104.340 58.035 105.340 ;
        RECT 56.705 103.890 57.165 104.150 ;
        RECT 56.305 103.345 56.565 103.665 ;
        RECT 57.305 103.595 57.535 104.340 ;
        RECT 58.200 104.150 58.430 105.545 ;
        RECT 58.685 105.340 58.915 105.345 ;
        RECT 58.595 104.340 58.915 105.340 ;
        RECT 59.095 105.340 59.325 105.935 ;
        RECT 59.465 105.545 59.925 105.775 ;
        RECT 59.095 104.340 59.415 105.340 ;
        RECT 58.085 103.890 58.545 104.150 ;
        RECT 56.705 103.365 57.535 103.595 ;
        RECT 56.335 103.160 56.565 103.345 ;
        RECT 56.335 102.160 56.655 103.160 ;
        RECT 54.800 96.895 56.050 99.975 ;
        RECT 56.335 99.630 56.565 102.160 ;
        RECT 56.820 102.000 57.050 103.365 ;
        RECT 57.685 103.345 57.945 103.665 ;
        RECT 58.685 103.595 58.915 104.340 ;
        RECT 59.580 104.150 59.810 105.545 ;
        RECT 60.065 105.340 60.295 105.345 ;
        RECT 59.975 104.340 60.295 105.340 ;
        RECT 60.475 105.340 60.705 105.935 ;
        RECT 60.845 105.545 61.305 105.775 ;
        RECT 60.475 104.340 60.795 105.340 ;
        RECT 59.465 103.890 59.925 104.150 ;
        RECT 58.085 103.365 58.915 103.595 ;
        RECT 57.305 103.160 57.535 103.165 ;
        RECT 57.215 102.160 57.535 103.160 ;
        RECT 56.705 101.680 57.165 102.000 ;
        RECT 56.705 99.775 57.165 100.035 ;
        RECT 56.335 98.980 56.655 99.630 ;
        RECT 56.820 98.820 57.050 99.775 ;
        RECT 57.305 99.630 57.535 102.160 ;
        RECT 57.215 98.980 57.535 99.630 ;
        RECT 57.715 103.160 57.945 103.345 ;
        RECT 57.715 102.160 58.035 103.160 ;
        RECT 57.715 99.630 57.945 102.160 ;
        RECT 58.200 102.000 58.430 103.365 ;
        RECT 59.065 103.345 59.325 103.665 ;
        RECT 60.065 103.595 60.295 104.340 ;
        RECT 60.960 104.150 61.190 105.545 ;
        RECT 61.445 105.340 61.675 105.345 ;
        RECT 61.355 104.340 61.675 105.340 ;
        RECT 61.855 105.340 62.085 105.935 ;
        RECT 62.225 105.545 62.685 105.775 ;
        RECT 61.855 104.340 62.175 105.340 ;
        RECT 60.845 103.890 61.305 104.150 ;
        RECT 59.465 103.365 60.295 103.595 ;
        RECT 58.685 103.160 58.915 103.165 ;
        RECT 58.595 102.160 58.915 103.160 ;
        RECT 58.085 101.680 58.545 102.000 ;
        RECT 58.085 99.775 58.545 100.035 ;
        RECT 57.715 98.980 58.035 99.630 ;
        RECT 58.200 98.820 58.430 99.775 ;
        RECT 58.685 99.630 58.915 102.160 ;
        RECT 58.595 98.980 58.915 99.630 ;
        RECT 59.095 103.160 59.325 103.345 ;
        RECT 59.095 102.160 59.415 103.160 ;
        RECT 59.095 99.630 59.325 102.160 ;
        RECT 59.580 102.000 59.810 103.365 ;
        RECT 60.445 103.345 60.705 103.665 ;
        RECT 61.445 103.595 61.675 104.340 ;
        RECT 62.340 104.150 62.570 105.545 ;
        RECT 62.825 105.340 63.055 105.345 ;
        RECT 62.735 104.340 63.055 105.340 ;
        RECT 63.235 105.340 63.465 105.935 ;
        RECT 63.605 105.545 64.065 105.775 ;
        RECT 63.235 104.340 63.555 105.340 ;
        RECT 62.225 103.890 62.685 104.150 ;
        RECT 60.845 103.365 61.675 103.595 ;
        RECT 60.065 103.160 60.295 103.165 ;
        RECT 59.975 102.160 60.295 103.160 ;
        RECT 59.465 101.680 59.925 102.000 ;
        RECT 59.465 99.775 59.925 100.035 ;
        RECT 59.095 98.980 59.415 99.630 ;
        RECT 59.580 98.820 59.810 99.775 ;
        RECT 60.065 99.630 60.295 102.160 ;
        RECT 59.975 98.980 60.295 99.630 ;
        RECT 60.475 103.160 60.705 103.345 ;
        RECT 60.475 102.160 60.795 103.160 ;
        RECT 60.475 99.630 60.705 102.160 ;
        RECT 60.960 102.000 61.190 103.365 ;
        RECT 61.825 103.345 62.085 103.665 ;
        RECT 62.825 103.595 63.055 104.340 ;
        RECT 63.720 104.150 63.950 105.545 ;
        RECT 64.205 105.340 64.435 105.345 ;
        RECT 64.115 104.340 64.435 105.340 ;
        RECT 64.615 105.340 64.845 105.935 ;
        RECT 64.985 105.545 65.445 105.775 ;
        RECT 64.615 104.340 64.935 105.340 ;
        RECT 63.605 103.890 64.065 104.150 ;
        RECT 62.225 103.365 63.055 103.595 ;
        RECT 61.445 103.160 61.675 103.165 ;
        RECT 61.355 102.160 61.675 103.160 ;
        RECT 60.845 101.680 61.305 102.000 ;
        RECT 60.845 99.775 61.305 100.035 ;
        RECT 60.475 98.980 60.795 99.630 ;
        RECT 60.960 98.820 61.190 99.775 ;
        RECT 61.445 99.630 61.675 102.160 ;
        RECT 61.355 98.980 61.675 99.630 ;
        RECT 61.855 103.160 62.085 103.345 ;
        RECT 61.855 102.160 62.175 103.160 ;
        RECT 61.855 99.630 62.085 102.160 ;
        RECT 62.340 102.000 62.570 103.365 ;
        RECT 63.205 103.345 63.465 103.665 ;
        RECT 64.205 103.595 64.435 104.340 ;
        RECT 65.100 104.150 65.330 105.545 ;
        RECT 65.585 105.340 65.815 105.345 ;
        RECT 65.495 104.340 65.815 105.340 ;
        RECT 65.995 105.340 66.225 105.935 ;
        RECT 66.365 105.545 66.825 105.775 ;
        RECT 65.995 104.340 66.315 105.340 ;
        RECT 64.985 103.890 65.445 104.150 ;
        RECT 63.605 103.365 64.435 103.595 ;
        RECT 62.825 103.160 63.055 103.165 ;
        RECT 62.735 102.160 63.055 103.160 ;
        RECT 62.225 101.680 62.685 102.000 ;
        RECT 62.225 99.775 62.685 100.035 ;
        RECT 61.855 98.980 62.175 99.630 ;
        RECT 62.340 98.820 62.570 99.775 ;
        RECT 62.825 99.630 63.055 102.160 ;
        RECT 62.735 98.980 63.055 99.630 ;
        RECT 63.235 103.160 63.465 103.345 ;
        RECT 63.235 102.160 63.555 103.160 ;
        RECT 63.235 99.630 63.465 102.160 ;
        RECT 63.720 102.000 63.950 103.365 ;
        RECT 64.585 103.345 64.845 103.665 ;
        RECT 65.585 103.595 65.815 104.340 ;
        RECT 66.480 104.150 66.710 105.545 ;
        RECT 66.965 105.340 67.195 105.345 ;
        RECT 66.875 104.340 67.195 105.340 ;
        RECT 67.375 105.340 67.605 105.935 ;
        RECT 67.745 105.545 68.205 105.775 ;
        RECT 67.375 104.340 67.695 105.340 ;
        RECT 66.365 103.890 66.825 104.150 ;
        RECT 64.985 103.365 65.815 103.595 ;
        RECT 64.205 103.160 64.435 103.165 ;
        RECT 64.115 102.160 64.435 103.160 ;
        RECT 63.605 101.680 64.065 102.000 ;
        RECT 63.605 99.775 64.065 100.035 ;
        RECT 63.235 98.980 63.555 99.630 ;
        RECT 63.720 98.820 63.950 99.775 ;
        RECT 64.205 99.630 64.435 102.160 ;
        RECT 64.115 98.980 64.435 99.630 ;
        RECT 64.615 103.160 64.845 103.345 ;
        RECT 64.615 102.160 64.935 103.160 ;
        RECT 64.615 99.630 64.845 102.160 ;
        RECT 65.100 102.000 65.330 103.365 ;
        RECT 65.965 103.345 66.225 103.665 ;
        RECT 66.965 103.595 67.195 104.340 ;
        RECT 67.860 104.150 68.090 105.545 ;
        RECT 68.345 105.340 68.575 105.345 ;
        RECT 68.255 104.340 68.575 105.340 ;
        RECT 68.755 105.340 68.985 105.935 ;
        RECT 69.125 105.545 69.585 105.775 ;
        RECT 68.755 104.340 69.075 105.340 ;
        RECT 67.745 103.890 68.205 104.150 ;
        RECT 66.365 103.365 67.195 103.595 ;
        RECT 65.585 103.160 65.815 103.165 ;
        RECT 65.495 102.160 65.815 103.160 ;
        RECT 64.985 101.680 65.445 102.000 ;
        RECT 64.985 99.775 65.445 100.035 ;
        RECT 64.615 98.980 64.935 99.630 ;
        RECT 65.100 98.820 65.330 99.775 ;
        RECT 65.585 99.630 65.815 102.160 ;
        RECT 65.495 98.980 65.815 99.630 ;
        RECT 65.995 103.160 66.225 103.345 ;
        RECT 65.995 102.160 66.315 103.160 ;
        RECT 65.995 99.630 66.225 102.160 ;
        RECT 66.480 102.000 66.710 103.365 ;
        RECT 67.345 103.345 67.605 103.665 ;
        RECT 68.345 103.595 68.575 104.340 ;
        RECT 69.240 104.150 69.470 105.545 ;
        RECT 69.725 105.340 69.955 105.345 ;
        RECT 69.635 104.340 69.955 105.340 ;
        RECT 70.135 105.340 70.365 105.935 ;
        RECT 70.505 105.545 70.965 105.775 ;
        RECT 70.135 104.340 70.455 105.340 ;
        RECT 69.125 103.890 69.585 104.150 ;
        RECT 67.745 103.365 68.575 103.595 ;
        RECT 66.965 103.160 67.195 103.165 ;
        RECT 66.875 102.160 67.195 103.160 ;
        RECT 66.365 101.680 66.825 102.000 ;
        RECT 66.365 99.775 66.825 100.035 ;
        RECT 65.995 98.980 66.315 99.630 ;
        RECT 66.480 98.820 66.710 99.775 ;
        RECT 66.965 99.630 67.195 102.160 ;
        RECT 66.875 98.980 67.195 99.630 ;
        RECT 67.375 103.160 67.605 103.345 ;
        RECT 67.375 102.160 67.695 103.160 ;
        RECT 67.375 99.630 67.605 102.160 ;
        RECT 67.860 102.000 68.090 103.365 ;
        RECT 68.725 103.345 68.985 103.665 ;
        RECT 69.725 103.595 69.955 104.340 ;
        RECT 70.620 104.150 70.850 105.545 ;
        RECT 71.105 105.340 71.335 105.345 ;
        RECT 71.015 104.340 71.335 105.340 ;
        RECT 71.515 105.340 71.745 105.935 ;
        RECT 71.885 105.545 72.345 105.775 ;
        RECT 71.515 104.340 71.835 105.340 ;
        RECT 70.505 103.890 70.965 104.150 ;
        RECT 69.125 103.365 69.955 103.595 ;
        RECT 68.345 103.160 68.575 103.165 ;
        RECT 68.255 102.160 68.575 103.160 ;
        RECT 67.745 101.680 68.205 102.000 ;
        RECT 67.745 99.775 68.205 100.035 ;
        RECT 67.375 98.980 67.695 99.630 ;
        RECT 67.860 98.820 68.090 99.775 ;
        RECT 68.345 99.630 68.575 102.160 ;
        RECT 68.255 98.980 68.575 99.630 ;
        RECT 68.755 103.160 68.985 103.345 ;
        RECT 68.755 102.160 69.075 103.160 ;
        RECT 68.755 99.630 68.985 102.160 ;
        RECT 69.240 102.000 69.470 103.365 ;
        RECT 70.105 103.345 70.365 103.665 ;
        RECT 71.105 103.595 71.335 104.340 ;
        RECT 72.000 104.150 72.230 105.545 ;
        RECT 72.485 105.340 72.715 105.345 ;
        RECT 72.395 104.340 72.715 105.340 ;
        RECT 72.895 105.340 73.125 105.935 ;
        RECT 73.265 105.545 73.725 105.775 ;
        RECT 72.895 104.340 73.215 105.340 ;
        RECT 71.885 103.890 72.345 104.150 ;
        RECT 70.505 103.365 71.335 103.595 ;
        RECT 69.725 103.160 69.955 103.165 ;
        RECT 69.635 102.160 69.955 103.160 ;
        RECT 69.125 101.680 69.585 102.000 ;
        RECT 69.125 99.775 69.585 100.035 ;
        RECT 68.755 98.980 69.075 99.630 ;
        RECT 69.240 98.820 69.470 99.775 ;
        RECT 69.725 99.630 69.955 102.160 ;
        RECT 69.635 98.980 69.955 99.630 ;
        RECT 70.135 103.160 70.365 103.345 ;
        RECT 70.135 102.160 70.455 103.160 ;
        RECT 70.135 99.630 70.365 102.160 ;
        RECT 70.620 102.000 70.850 103.365 ;
        RECT 71.485 103.345 71.745 103.665 ;
        RECT 72.485 103.595 72.715 104.340 ;
        RECT 73.380 104.150 73.610 105.545 ;
        RECT 73.865 105.340 74.095 105.345 ;
        RECT 73.775 104.340 74.095 105.340 ;
        RECT 74.275 105.340 74.505 105.935 ;
        RECT 74.645 105.545 75.105 105.775 ;
        RECT 74.275 104.340 74.595 105.340 ;
        RECT 73.265 103.890 73.725 104.150 ;
        RECT 71.885 103.365 72.715 103.595 ;
        RECT 71.105 103.160 71.335 103.165 ;
        RECT 71.015 102.160 71.335 103.160 ;
        RECT 70.505 101.680 70.965 102.000 ;
        RECT 70.505 99.775 70.965 100.035 ;
        RECT 70.135 98.980 70.455 99.630 ;
        RECT 70.620 98.820 70.850 99.775 ;
        RECT 71.105 99.630 71.335 102.160 ;
        RECT 71.015 98.980 71.335 99.630 ;
        RECT 71.515 103.160 71.745 103.345 ;
        RECT 71.515 102.160 71.835 103.160 ;
        RECT 71.515 99.630 71.745 102.160 ;
        RECT 72.000 102.000 72.230 103.365 ;
        RECT 72.865 103.345 73.125 103.665 ;
        RECT 73.865 103.595 74.095 104.340 ;
        RECT 74.760 104.150 74.990 105.545 ;
        RECT 75.245 105.340 75.475 105.345 ;
        RECT 75.155 104.340 75.475 105.340 ;
        RECT 75.655 105.340 75.885 105.935 ;
        RECT 76.025 105.545 76.485 105.775 ;
        RECT 75.655 104.340 75.975 105.340 ;
        RECT 74.645 103.890 75.105 104.150 ;
        RECT 73.265 103.365 74.095 103.595 ;
        RECT 72.485 103.160 72.715 103.165 ;
        RECT 72.395 102.160 72.715 103.160 ;
        RECT 71.885 101.680 72.345 102.000 ;
        RECT 71.885 99.775 72.345 100.035 ;
        RECT 71.515 98.980 71.835 99.630 ;
        RECT 72.000 98.820 72.230 99.775 ;
        RECT 72.485 99.630 72.715 102.160 ;
        RECT 72.395 98.980 72.715 99.630 ;
        RECT 72.895 103.160 73.125 103.345 ;
        RECT 72.895 102.160 73.215 103.160 ;
        RECT 72.895 99.630 73.125 102.160 ;
        RECT 73.380 102.000 73.610 103.365 ;
        RECT 74.245 103.345 74.505 103.665 ;
        RECT 75.245 103.595 75.475 104.340 ;
        RECT 76.140 104.150 76.370 105.545 ;
        RECT 76.625 105.340 76.855 105.345 ;
        RECT 76.535 104.340 76.855 105.340 ;
        RECT 77.035 105.340 77.265 105.935 ;
        RECT 77.405 105.545 77.865 105.775 ;
        RECT 77.035 104.340 77.355 105.340 ;
        RECT 76.025 103.890 76.485 104.150 ;
        RECT 74.645 103.365 75.475 103.595 ;
        RECT 73.865 103.160 74.095 103.165 ;
        RECT 73.775 102.160 74.095 103.160 ;
        RECT 73.265 101.680 73.725 102.000 ;
        RECT 73.265 99.775 73.725 100.035 ;
        RECT 72.895 98.980 73.215 99.630 ;
        RECT 73.380 98.820 73.610 99.775 ;
        RECT 73.865 99.630 74.095 102.160 ;
        RECT 73.775 98.980 74.095 99.630 ;
        RECT 74.275 103.160 74.505 103.345 ;
        RECT 74.275 102.160 74.595 103.160 ;
        RECT 74.275 99.630 74.505 102.160 ;
        RECT 74.760 102.000 74.990 103.365 ;
        RECT 75.625 103.345 75.885 103.665 ;
        RECT 76.625 103.595 76.855 104.340 ;
        RECT 77.520 104.150 77.750 105.545 ;
        RECT 78.005 105.340 78.235 105.345 ;
        RECT 77.915 104.340 78.235 105.340 ;
        RECT 78.415 105.340 78.645 105.935 ;
        RECT 78.785 105.545 79.245 105.775 ;
        RECT 78.415 104.340 78.735 105.340 ;
        RECT 77.405 103.890 77.865 104.150 ;
        RECT 76.025 103.365 76.855 103.595 ;
        RECT 75.245 103.160 75.475 103.165 ;
        RECT 75.155 102.160 75.475 103.160 ;
        RECT 74.645 101.680 75.105 102.000 ;
        RECT 74.645 99.775 75.105 100.035 ;
        RECT 74.275 98.980 74.595 99.630 ;
        RECT 74.760 98.820 74.990 99.775 ;
        RECT 75.245 99.630 75.475 102.160 ;
        RECT 75.155 98.980 75.475 99.630 ;
        RECT 75.655 103.160 75.885 103.345 ;
        RECT 75.655 102.160 75.975 103.160 ;
        RECT 75.655 99.630 75.885 102.160 ;
        RECT 76.140 102.000 76.370 103.365 ;
        RECT 77.005 103.345 77.265 103.665 ;
        RECT 78.005 103.595 78.235 104.340 ;
        RECT 78.900 104.150 79.130 105.545 ;
        RECT 79.385 105.340 79.615 105.345 ;
        RECT 79.295 104.340 79.615 105.340 ;
        RECT 79.795 105.340 80.025 105.935 ;
        RECT 80.165 105.545 80.625 105.775 ;
        RECT 79.795 104.340 80.115 105.340 ;
        RECT 78.785 103.890 79.245 104.150 ;
        RECT 77.405 103.365 78.235 103.595 ;
        RECT 76.625 103.160 76.855 103.165 ;
        RECT 76.535 102.160 76.855 103.160 ;
        RECT 76.025 101.680 76.485 102.000 ;
        RECT 76.025 99.775 76.485 100.035 ;
        RECT 75.655 98.980 75.975 99.630 ;
        RECT 76.140 98.820 76.370 99.775 ;
        RECT 76.625 99.630 76.855 102.160 ;
        RECT 76.535 98.980 76.855 99.630 ;
        RECT 77.035 103.160 77.265 103.345 ;
        RECT 77.035 102.160 77.355 103.160 ;
        RECT 77.035 99.630 77.265 102.160 ;
        RECT 77.520 102.000 77.750 103.365 ;
        RECT 78.385 103.345 78.645 103.665 ;
        RECT 79.385 103.595 79.615 104.340 ;
        RECT 80.280 104.150 80.510 105.545 ;
        RECT 80.765 105.340 80.995 105.345 ;
        RECT 80.675 104.340 80.995 105.340 ;
        RECT 81.175 105.340 81.405 105.935 ;
        RECT 81.545 105.545 82.005 105.775 ;
        RECT 81.175 104.340 81.495 105.340 ;
        RECT 80.165 103.890 80.625 104.150 ;
        RECT 78.785 103.365 79.615 103.595 ;
        RECT 78.005 103.160 78.235 103.165 ;
        RECT 77.915 102.160 78.235 103.160 ;
        RECT 77.405 101.680 77.865 102.000 ;
        RECT 77.405 99.775 77.865 100.035 ;
        RECT 77.035 98.980 77.355 99.630 ;
        RECT 77.520 98.820 77.750 99.775 ;
        RECT 78.005 99.630 78.235 102.160 ;
        RECT 77.915 98.980 78.235 99.630 ;
        RECT 78.415 103.160 78.645 103.345 ;
        RECT 78.415 102.160 78.735 103.160 ;
        RECT 78.415 99.630 78.645 102.160 ;
        RECT 78.900 102.000 79.130 103.365 ;
        RECT 79.765 103.345 80.025 103.665 ;
        RECT 80.765 103.595 80.995 104.340 ;
        RECT 81.660 104.150 81.890 105.545 ;
        RECT 82.145 105.340 82.375 105.345 ;
        RECT 82.055 104.340 82.375 105.340 ;
        RECT 81.545 103.890 82.005 104.150 ;
        RECT 80.165 103.365 80.995 103.595 ;
        RECT 79.385 103.160 79.615 103.165 ;
        RECT 79.295 102.160 79.615 103.160 ;
        RECT 78.785 101.680 79.245 102.000 ;
        RECT 78.785 99.775 79.245 100.035 ;
        RECT 78.415 98.980 78.735 99.630 ;
        RECT 78.900 98.820 79.130 99.775 ;
        RECT 79.385 99.630 79.615 102.160 ;
        RECT 79.295 98.980 79.615 99.630 ;
        RECT 79.795 103.160 80.025 103.345 ;
        RECT 79.795 102.160 80.115 103.160 ;
        RECT 79.795 99.630 80.025 102.160 ;
        RECT 80.280 102.000 80.510 103.365 ;
        RECT 81.145 103.345 81.405 103.665 ;
        RECT 82.145 103.595 82.375 104.340 ;
        RECT 81.545 103.365 82.375 103.595 ;
        RECT 80.765 103.160 80.995 103.165 ;
        RECT 80.675 102.160 80.995 103.160 ;
        RECT 80.165 101.680 80.625 102.000 ;
        RECT 80.165 99.775 80.625 100.035 ;
        RECT 79.795 98.980 80.115 99.630 ;
        RECT 80.280 98.820 80.510 99.775 ;
        RECT 80.765 99.630 80.995 102.160 ;
        RECT 80.675 98.980 80.995 99.630 ;
        RECT 81.175 103.160 81.405 103.345 ;
        RECT 81.175 102.160 81.495 103.160 ;
        RECT 81.175 99.630 81.405 102.160 ;
        RECT 81.660 102.000 81.890 103.365 ;
        RECT 82.145 103.160 82.375 103.165 ;
        RECT 82.055 102.160 82.375 103.160 ;
        RECT 81.545 101.680 82.005 102.000 ;
        RECT 81.545 99.775 82.005 100.035 ;
        RECT 81.175 98.980 81.495 99.630 ;
        RECT 81.660 98.820 81.890 99.775 ;
        RECT 82.145 99.630 82.375 102.160 ;
        RECT 82.660 101.815 83.160 106.140 ;
        RECT 82.055 98.980 82.375 99.630 ;
        RECT 56.705 98.590 57.165 98.820 ;
        RECT 58.085 98.590 58.545 98.820 ;
        RECT 59.465 98.590 59.925 98.820 ;
        RECT 60.845 98.590 61.305 98.820 ;
        RECT 62.225 98.590 62.685 98.820 ;
        RECT 63.605 98.590 64.065 98.820 ;
        RECT 64.985 98.590 65.445 98.820 ;
        RECT 66.365 98.590 66.825 98.820 ;
        RECT 67.745 98.590 68.205 98.820 ;
        RECT 69.125 98.590 69.585 98.820 ;
        RECT 70.505 98.590 70.965 98.820 ;
        RECT 71.885 98.590 72.345 98.820 ;
        RECT 73.265 98.590 73.725 98.820 ;
        RECT 74.645 98.590 75.105 98.820 ;
        RECT 76.025 98.590 76.485 98.820 ;
        RECT 77.405 98.590 77.865 98.820 ;
        RECT 78.785 98.590 79.245 98.820 ;
        RECT 80.165 98.590 80.625 98.820 ;
        RECT 81.545 98.590 82.005 98.820 ;
        RECT 56.705 98.280 57.050 98.590 ;
        RECT 58.085 98.280 58.430 98.590 ;
        RECT 59.465 98.280 59.810 98.590 ;
        RECT 60.845 98.280 61.190 98.590 ;
        RECT 62.225 98.280 62.570 98.590 ;
        RECT 63.605 98.280 63.950 98.590 ;
        RECT 64.985 98.280 65.330 98.590 ;
        RECT 66.365 98.280 66.710 98.590 ;
        RECT 67.745 98.280 68.090 98.590 ;
        RECT 69.125 98.280 69.470 98.590 ;
        RECT 70.505 98.280 70.850 98.590 ;
        RECT 71.885 98.280 72.230 98.590 ;
        RECT 73.265 98.280 73.610 98.590 ;
        RECT 74.645 98.280 74.990 98.590 ;
        RECT 76.025 98.280 76.370 98.590 ;
        RECT 77.405 98.280 77.750 98.590 ;
        RECT 78.785 98.280 79.130 98.590 ;
        RECT 80.165 98.280 80.510 98.590 ;
        RECT 81.545 98.280 81.890 98.590 ;
        RECT 56.705 98.050 57.165 98.280 ;
        RECT 58.085 98.050 58.545 98.280 ;
        RECT 59.465 98.050 59.925 98.280 ;
        RECT 60.845 98.050 61.305 98.280 ;
        RECT 62.225 98.050 62.685 98.280 ;
        RECT 63.605 98.050 64.065 98.280 ;
        RECT 64.985 98.050 65.445 98.280 ;
        RECT 66.365 98.050 66.825 98.280 ;
        RECT 67.745 98.050 68.205 98.280 ;
        RECT 69.125 98.050 69.585 98.280 ;
        RECT 70.505 98.050 70.965 98.280 ;
        RECT 71.885 98.050 72.345 98.280 ;
        RECT 73.265 98.050 73.725 98.280 ;
        RECT 74.645 98.050 75.105 98.280 ;
        RECT 76.025 98.050 76.485 98.280 ;
        RECT 77.405 98.050 77.865 98.280 ;
        RECT 78.785 98.050 79.245 98.280 ;
        RECT 80.165 98.050 80.625 98.280 ;
        RECT 81.545 98.050 82.005 98.280 ;
        RECT 56.335 97.240 56.655 97.890 ;
        RECT 56.335 96.645 56.565 97.240 ;
        RECT 56.820 97.080 57.050 98.050 ;
        RECT 57.215 97.240 57.535 97.890 ;
        RECT 57.715 97.240 58.035 97.890 ;
        RECT 56.705 96.850 57.165 97.080 ;
        RECT 57.715 96.645 57.945 97.240 ;
        RECT 58.200 97.080 58.430 98.050 ;
        RECT 58.595 97.240 58.915 97.890 ;
        RECT 59.095 97.240 59.415 97.890 ;
        RECT 58.085 96.850 58.545 97.080 ;
        RECT 59.095 96.645 59.325 97.240 ;
        RECT 59.580 97.080 59.810 98.050 ;
        RECT 59.975 97.240 60.295 97.890 ;
        RECT 60.475 97.240 60.795 97.890 ;
        RECT 59.465 96.850 59.925 97.080 ;
        RECT 60.475 96.645 60.705 97.240 ;
        RECT 60.960 97.080 61.190 98.050 ;
        RECT 61.355 97.240 61.675 97.890 ;
        RECT 61.855 97.240 62.175 97.890 ;
        RECT 60.845 96.850 61.305 97.080 ;
        RECT 61.855 96.645 62.085 97.240 ;
        RECT 62.340 97.080 62.570 98.050 ;
        RECT 62.735 97.240 63.055 97.890 ;
        RECT 63.235 97.240 63.555 97.890 ;
        RECT 62.225 96.850 62.685 97.080 ;
        RECT 63.235 96.645 63.465 97.240 ;
        RECT 63.720 97.080 63.950 98.050 ;
        RECT 64.115 97.240 64.435 97.890 ;
        RECT 64.615 97.240 64.935 97.890 ;
        RECT 63.605 96.850 64.065 97.080 ;
        RECT 64.615 96.645 64.845 97.240 ;
        RECT 65.100 97.080 65.330 98.050 ;
        RECT 65.495 97.240 65.815 97.890 ;
        RECT 65.995 97.240 66.315 97.890 ;
        RECT 64.985 96.850 65.445 97.080 ;
        RECT 65.995 96.645 66.225 97.240 ;
        RECT 66.480 97.080 66.710 98.050 ;
        RECT 66.875 97.240 67.195 97.890 ;
        RECT 67.375 97.240 67.695 97.890 ;
        RECT 66.365 96.850 66.825 97.080 ;
        RECT 67.375 96.645 67.605 97.240 ;
        RECT 67.860 97.080 68.090 98.050 ;
        RECT 68.255 97.240 68.575 97.890 ;
        RECT 68.755 97.240 69.075 97.890 ;
        RECT 67.745 96.850 68.205 97.080 ;
        RECT 68.755 96.645 68.985 97.240 ;
        RECT 69.240 97.080 69.470 98.050 ;
        RECT 69.635 97.240 69.955 97.890 ;
        RECT 70.135 97.240 70.455 97.890 ;
        RECT 69.125 96.850 69.585 97.080 ;
        RECT 70.135 96.645 70.365 97.240 ;
        RECT 70.620 97.080 70.850 98.050 ;
        RECT 71.015 97.240 71.335 97.890 ;
        RECT 71.515 97.240 71.835 97.890 ;
        RECT 70.505 96.850 70.965 97.080 ;
        RECT 71.515 96.645 71.745 97.240 ;
        RECT 72.000 97.080 72.230 98.050 ;
        RECT 72.395 97.240 72.715 97.890 ;
        RECT 72.895 97.240 73.215 97.890 ;
        RECT 71.885 96.850 72.345 97.080 ;
        RECT 72.895 96.645 73.125 97.240 ;
        RECT 73.380 97.080 73.610 98.050 ;
        RECT 73.775 97.240 74.095 97.890 ;
        RECT 74.275 97.240 74.595 97.890 ;
        RECT 73.265 96.850 73.725 97.080 ;
        RECT 74.275 96.645 74.505 97.240 ;
        RECT 74.760 97.080 74.990 98.050 ;
        RECT 75.155 97.240 75.475 97.890 ;
        RECT 75.655 97.240 75.975 97.890 ;
        RECT 74.645 96.850 75.105 97.080 ;
        RECT 75.655 96.645 75.885 97.240 ;
        RECT 76.140 97.080 76.370 98.050 ;
        RECT 76.535 97.240 76.855 97.890 ;
        RECT 77.035 97.240 77.355 97.890 ;
        RECT 76.025 96.850 76.485 97.080 ;
        RECT 77.035 96.645 77.265 97.240 ;
        RECT 77.520 97.080 77.750 98.050 ;
        RECT 77.915 97.240 78.235 97.890 ;
        RECT 78.415 97.240 78.735 97.890 ;
        RECT 77.405 96.850 77.865 97.080 ;
        RECT 78.415 96.645 78.645 97.240 ;
        RECT 78.900 97.080 79.130 98.050 ;
        RECT 79.295 97.240 79.615 97.890 ;
        RECT 79.795 97.240 80.115 97.890 ;
        RECT 78.785 96.850 79.245 97.080 ;
        RECT 79.795 96.645 80.025 97.240 ;
        RECT 80.280 97.080 80.510 98.050 ;
        RECT 80.675 97.240 80.995 97.890 ;
        RECT 81.175 97.240 81.495 97.890 ;
        RECT 80.165 96.850 80.625 97.080 ;
        RECT 81.175 96.645 81.405 97.240 ;
        RECT 81.660 97.080 81.890 98.050 ;
        RECT 82.055 97.240 82.375 97.890 ;
        RECT 81.545 96.850 82.005 97.080 ;
        RECT 82.660 96.895 83.910 99.975 ;
        RECT 56.245 96.355 82.465 96.645 ;
        RECT 68.970 95.390 69.230 95.465 ;
        RECT 71.140 95.390 71.400 95.465 ;
        RECT 68.970 95.220 71.400 95.390 ;
        RECT 68.970 95.145 69.230 95.220 ;
        RECT 71.140 95.145 71.400 95.220 ;
        RECT 35.140 95.005 35.400 95.080 ;
        RECT 57.930 95.005 58.190 95.080 ;
        RECT 35.140 94.835 58.190 95.005 ;
        RECT 35.140 94.760 35.400 94.835 ;
        RECT 57.930 94.760 58.190 94.835 ;
        RECT 70.350 95.005 70.610 95.080 ;
        RECT 75.255 95.005 75.515 95.080 ;
        RECT 70.350 94.835 75.515 95.005 ;
        RECT 70.350 94.760 70.610 94.835 ;
        RECT 75.255 94.760 75.515 94.835 ;
        RECT 39.640 94.620 39.900 94.695 ;
        RECT 59.310 94.620 59.570 94.695 ;
        RECT 39.640 94.450 59.570 94.620 ;
        RECT 39.640 94.375 39.900 94.450 ;
        RECT 59.310 94.375 59.570 94.450 ;
        RECT 71.730 94.620 71.990 94.695 ;
        RECT 80.525 94.620 80.785 94.695 ;
        RECT 71.730 94.450 80.785 94.620 ;
        RECT 71.730 94.375 71.990 94.450 ;
        RECT 80.525 94.375 80.785 94.450 ;
        RECT 44.140 94.235 44.400 94.310 ;
        RECT 60.690 94.235 60.950 94.310 ;
        RECT 44.140 94.065 60.950 94.235 ;
        RECT 44.140 93.990 44.400 94.065 ;
        RECT 60.690 93.990 60.950 94.065 ;
        RECT 73.110 94.235 73.370 94.310 ;
        RECT 84.640 94.235 84.900 94.310 ;
        RECT 73.110 94.065 84.900 94.235 ;
        RECT 73.110 93.990 73.370 94.065 ;
        RECT 84.640 93.990 84.900 94.065 ;
        RECT 48.640 93.850 48.900 93.925 ;
        RECT 62.070 93.850 62.330 93.925 ;
        RECT 48.640 93.680 62.330 93.850 ;
        RECT 48.640 93.605 48.900 93.680 ;
        RECT 62.070 93.605 62.330 93.680 ;
        RECT 74.490 93.850 74.750 93.925 ;
        RECT 89.140 93.850 89.400 93.925 ;
        RECT 74.490 93.680 89.400 93.850 ;
        RECT 74.490 93.605 74.750 93.680 ;
        RECT 89.140 93.605 89.400 93.680 ;
        RECT 53.140 93.465 53.400 93.540 ;
        RECT 63.450 93.465 63.710 93.540 ;
        RECT 53.140 93.295 63.710 93.465 ;
        RECT 53.140 93.220 53.400 93.295 ;
        RECT 63.450 93.220 63.710 93.295 ;
        RECT 75.870 93.465 76.130 93.540 ;
        RECT 93.640 93.465 93.900 93.540 ;
        RECT 75.870 93.295 93.900 93.465 ;
        RECT 75.870 93.220 76.130 93.295 ;
        RECT 93.640 93.220 93.900 93.295 ;
        RECT 57.640 93.080 57.900 93.155 ;
        RECT 64.830 93.080 65.090 93.155 ;
        RECT 57.640 92.910 65.090 93.080 ;
        RECT 57.640 92.835 57.900 92.910 ;
        RECT 64.830 92.835 65.090 92.910 ;
        RECT 77.250 93.080 77.510 93.155 ;
        RECT 98.140 93.080 98.400 93.155 ;
        RECT 77.250 92.910 98.400 93.080 ;
        RECT 77.250 92.835 77.510 92.910 ;
        RECT 98.140 92.835 98.400 92.910 ;
        RECT 62.140 92.695 62.400 92.770 ;
        RECT 66.210 92.695 66.470 92.770 ;
        RECT 62.140 92.525 66.470 92.695 ;
        RECT 62.140 92.450 62.400 92.525 ;
        RECT 66.210 92.450 66.470 92.525 ;
        RECT 78.630 92.695 78.890 92.770 ;
        RECT 102.640 92.695 102.900 92.770 ;
        RECT 78.630 92.525 102.900 92.695 ;
        RECT 78.630 92.450 78.890 92.525 ;
        RECT 102.640 92.450 102.900 92.525 ;
        RECT 66.640 92.310 66.900 92.385 ;
        RECT 67.590 92.310 67.850 92.385 ;
        RECT 66.640 92.140 67.850 92.310 ;
        RECT 66.640 92.065 66.900 92.140 ;
        RECT 67.590 92.065 67.850 92.140 ;
        RECT 80.010 92.310 80.270 92.385 ;
        RECT 107.140 92.310 107.400 92.385 ;
        RECT 80.010 92.140 107.400 92.310 ;
        RECT 80.010 92.065 80.270 92.140 ;
        RECT 107.140 92.065 107.400 92.140 ;
        RECT 31.065 91.455 107.565 91.745 ;
        RECT 30.640 89.440 30.960 91.280 ;
        RECT 31.275 90.860 31.445 91.455 ;
        RECT 31.585 91.065 32.045 91.295 ;
        RECT 33.085 91.065 33.545 91.295 ;
        RECT 31.245 89.860 31.475 90.860 ;
        RECT 31.275 89.840 31.445 89.860 ;
        RECT 31.730 89.655 31.900 91.065 ;
        RECT 32.185 90.860 32.355 90.880 ;
        RECT 32.775 90.860 32.945 90.880 ;
        RECT 32.155 90.445 32.385 90.860 ;
        RECT 32.745 90.445 32.975 90.860 ;
        RECT 32.155 90.275 32.975 90.445 ;
        RECT 32.155 89.860 32.385 90.275 ;
        RECT 32.745 89.860 32.975 90.275 ;
        RECT 32.185 89.840 32.355 89.860 ;
        RECT 32.775 89.840 32.945 89.860 ;
        RECT 33.230 89.655 33.400 91.065 ;
        RECT 33.685 90.860 33.855 90.880 ;
        RECT 34.275 90.860 34.445 91.455 ;
        RECT 34.585 91.065 35.045 91.295 ;
        RECT 33.655 89.860 33.885 90.860 ;
        RECT 34.245 89.860 34.475 90.860 ;
        RECT 31.585 89.425 32.045 89.655 ;
        RECT 33.085 89.425 33.545 89.655 ;
        RECT 30.550 84.695 30.850 87.740 ;
        RECT 31.730 87.720 31.900 89.425 ;
        RECT 32.110 88.465 32.430 88.725 ;
        RECT 31.585 87.490 32.045 87.720 ;
        RECT 31.275 87.330 31.445 87.350 ;
        RECT 31.245 86.680 31.475 87.330 ;
        RECT 31.275 86.085 31.445 86.680 ;
        RECT 31.730 86.565 31.900 87.490 ;
        RECT 32.185 87.330 32.355 88.465 ;
        RECT 33.230 87.720 33.400 89.425 ;
        RECT 33.685 88.725 33.855 89.860 ;
        RECT 34.275 89.840 34.445 89.860 ;
        RECT 34.730 89.655 34.900 91.065 ;
        RECT 35.140 90.635 35.400 90.955 ;
        RECT 35.775 90.860 35.945 91.455 ;
        RECT 36.085 91.065 36.545 91.295 ;
        RECT 37.585 91.065 38.045 91.295 ;
        RECT 35.155 89.860 35.385 90.635 ;
        RECT 35.745 89.860 35.975 90.860 ;
        RECT 34.585 89.425 35.045 89.655 ;
        RECT 34.730 88.725 34.900 89.425 ;
        RECT 33.610 88.465 33.930 88.725 ;
        RECT 34.655 88.465 34.975 88.725 ;
        RECT 33.085 87.490 33.545 87.720 ;
        RECT 32.775 87.330 32.945 87.350 ;
        RECT 32.155 86.680 32.385 87.330 ;
        RECT 32.745 86.680 32.975 87.330 ;
        RECT 32.185 86.660 32.355 86.680 ;
        RECT 31.685 86.520 31.945 86.565 ;
        RECT 31.585 86.290 32.045 86.520 ;
        RECT 31.685 86.245 31.945 86.290 ;
        RECT 31.685 86.085 31.945 86.100 ;
        RECT 32.775 86.085 32.945 86.680 ;
        RECT 33.230 86.565 33.400 87.490 ;
        RECT 33.685 87.330 33.855 88.465 ;
        RECT 34.730 87.720 34.900 88.465 ;
        RECT 34.585 87.490 35.045 87.720 ;
        RECT 34.275 87.330 34.445 87.350 ;
        RECT 33.655 86.680 33.885 87.330 ;
        RECT 34.245 86.680 34.475 87.330 ;
        RECT 33.685 86.660 33.855 86.680 ;
        RECT 33.185 86.520 33.445 86.565 ;
        RECT 33.085 86.290 33.545 86.520 ;
        RECT 33.185 86.245 33.445 86.290 ;
        RECT 34.275 86.085 34.445 86.680 ;
        RECT 34.730 86.520 34.900 87.490 ;
        RECT 35.185 87.330 35.355 89.860 ;
        RECT 35.775 89.840 35.945 89.860 ;
        RECT 36.230 89.655 36.400 91.065 ;
        RECT 36.685 90.860 36.855 90.880 ;
        RECT 37.275 90.860 37.445 90.880 ;
        RECT 36.655 90.445 36.885 90.860 ;
        RECT 37.245 90.445 37.475 90.860 ;
        RECT 36.655 90.275 37.475 90.445 ;
        RECT 36.655 89.860 36.885 90.275 ;
        RECT 37.245 89.860 37.475 90.275 ;
        RECT 36.685 89.840 36.855 89.860 ;
        RECT 37.275 89.840 37.445 89.860 ;
        RECT 37.730 89.655 37.900 91.065 ;
        RECT 38.185 90.860 38.355 90.880 ;
        RECT 38.775 90.860 38.945 91.455 ;
        RECT 39.085 91.065 39.545 91.295 ;
        RECT 38.155 89.860 38.385 90.860 ;
        RECT 38.745 89.860 38.975 90.860 ;
        RECT 36.085 89.425 36.545 89.655 ;
        RECT 37.585 89.425 38.045 89.655 ;
        RECT 36.230 87.720 36.400 89.425 ;
        RECT 36.610 88.465 36.930 88.725 ;
        RECT 36.085 87.490 36.545 87.720 ;
        RECT 35.775 87.330 35.945 87.350 ;
        RECT 35.155 86.680 35.385 87.330 ;
        RECT 35.745 86.680 35.975 87.330 ;
        RECT 35.185 86.660 35.355 86.680 ;
        RECT 34.585 86.290 35.045 86.520 ;
        RECT 35.775 86.085 35.945 86.680 ;
        RECT 36.230 86.565 36.400 87.490 ;
        RECT 36.685 87.330 36.855 88.465 ;
        RECT 37.730 87.720 37.900 89.425 ;
        RECT 38.185 88.725 38.355 89.860 ;
        RECT 38.775 89.840 38.945 89.860 ;
        RECT 39.230 89.655 39.400 91.065 ;
        RECT 39.640 90.635 39.900 90.955 ;
        RECT 40.275 90.860 40.445 91.455 ;
        RECT 40.585 91.065 41.045 91.295 ;
        RECT 42.085 91.065 42.545 91.295 ;
        RECT 39.655 89.860 39.885 90.635 ;
        RECT 40.245 89.860 40.475 90.860 ;
        RECT 39.085 89.425 39.545 89.655 ;
        RECT 39.230 88.725 39.400 89.425 ;
        RECT 38.110 88.465 38.430 88.725 ;
        RECT 39.155 88.465 39.475 88.725 ;
        RECT 37.585 87.490 38.045 87.720 ;
        RECT 37.275 87.330 37.445 87.350 ;
        RECT 36.655 86.680 36.885 87.330 ;
        RECT 37.245 86.680 37.475 87.330 ;
        RECT 36.685 86.660 36.855 86.680 ;
        RECT 36.185 86.520 36.445 86.565 ;
        RECT 36.085 86.290 36.545 86.520 ;
        RECT 36.185 86.245 36.445 86.290 ;
        RECT 37.275 86.085 37.445 86.680 ;
        RECT 37.730 86.565 37.900 87.490 ;
        RECT 38.185 87.330 38.355 88.465 ;
        RECT 39.230 87.720 39.400 88.465 ;
        RECT 39.085 87.490 39.545 87.720 ;
        RECT 38.775 87.330 38.945 87.350 ;
        RECT 38.155 86.680 38.385 87.330 ;
        RECT 38.745 86.680 38.975 87.330 ;
        RECT 38.185 86.660 38.355 86.680 ;
        RECT 37.685 86.520 37.945 86.565 ;
        RECT 37.585 86.290 38.045 86.520 ;
        RECT 37.685 86.245 37.945 86.290 ;
        RECT 38.775 86.085 38.945 86.680 ;
        RECT 39.230 86.520 39.400 87.490 ;
        RECT 39.685 87.330 39.855 89.860 ;
        RECT 40.275 89.840 40.445 89.860 ;
        RECT 40.730 89.655 40.900 91.065 ;
        RECT 41.185 90.860 41.355 90.880 ;
        RECT 41.775 90.860 41.945 90.880 ;
        RECT 41.155 90.445 41.385 90.860 ;
        RECT 41.745 90.445 41.975 90.860 ;
        RECT 41.155 90.275 41.975 90.445 ;
        RECT 41.155 89.860 41.385 90.275 ;
        RECT 41.745 89.860 41.975 90.275 ;
        RECT 41.185 89.840 41.355 89.860 ;
        RECT 41.775 89.840 41.945 89.860 ;
        RECT 42.230 89.655 42.400 91.065 ;
        RECT 42.685 90.860 42.855 90.880 ;
        RECT 43.275 90.860 43.445 91.455 ;
        RECT 43.585 91.065 44.045 91.295 ;
        RECT 42.655 89.860 42.885 90.860 ;
        RECT 43.245 89.860 43.475 90.860 ;
        RECT 40.585 89.425 41.045 89.655 ;
        RECT 42.085 89.425 42.545 89.655 ;
        RECT 40.730 87.720 40.900 89.425 ;
        RECT 41.110 88.465 41.430 88.725 ;
        RECT 40.585 87.490 41.045 87.720 ;
        RECT 40.275 87.330 40.445 87.350 ;
        RECT 39.655 86.680 39.885 87.330 ;
        RECT 40.245 86.680 40.475 87.330 ;
        RECT 39.685 86.660 39.855 86.680 ;
        RECT 39.085 86.290 39.545 86.520 ;
        RECT 40.275 86.085 40.445 86.680 ;
        RECT 40.730 86.565 40.900 87.490 ;
        RECT 41.185 87.330 41.355 88.465 ;
        RECT 42.230 87.720 42.400 89.425 ;
        RECT 42.685 88.725 42.855 89.860 ;
        RECT 43.275 89.840 43.445 89.860 ;
        RECT 43.730 89.655 43.900 91.065 ;
        RECT 44.140 90.635 44.400 90.955 ;
        RECT 44.775 90.860 44.945 91.455 ;
        RECT 45.085 91.065 45.545 91.295 ;
        RECT 46.585 91.065 47.045 91.295 ;
        RECT 44.155 89.860 44.385 90.635 ;
        RECT 44.745 89.860 44.975 90.860 ;
        RECT 43.585 89.425 44.045 89.655 ;
        RECT 43.730 88.725 43.900 89.425 ;
        RECT 42.610 88.465 42.930 88.725 ;
        RECT 43.655 88.465 43.975 88.725 ;
        RECT 42.085 87.490 42.545 87.720 ;
        RECT 41.775 87.330 41.945 87.350 ;
        RECT 41.155 86.680 41.385 87.330 ;
        RECT 41.745 86.680 41.975 87.330 ;
        RECT 41.185 86.660 41.355 86.680 ;
        RECT 40.685 86.520 40.945 86.565 ;
        RECT 40.585 86.290 41.045 86.520 ;
        RECT 40.685 86.245 40.945 86.290 ;
        RECT 41.775 86.085 41.945 86.680 ;
        RECT 42.230 86.565 42.400 87.490 ;
        RECT 42.685 87.330 42.855 88.465 ;
        RECT 43.730 87.720 43.900 88.465 ;
        RECT 43.585 87.490 44.045 87.720 ;
        RECT 43.275 87.330 43.445 87.350 ;
        RECT 42.655 86.680 42.885 87.330 ;
        RECT 43.245 86.680 43.475 87.330 ;
        RECT 42.685 86.660 42.855 86.680 ;
        RECT 42.185 86.520 42.445 86.565 ;
        RECT 42.085 86.290 42.545 86.520 ;
        RECT 42.185 86.245 42.445 86.290 ;
        RECT 43.275 86.085 43.445 86.680 ;
        RECT 43.730 86.520 43.900 87.490 ;
        RECT 44.185 87.330 44.355 89.860 ;
        RECT 44.775 89.840 44.945 89.860 ;
        RECT 45.230 89.655 45.400 91.065 ;
        RECT 45.685 90.860 45.855 90.880 ;
        RECT 46.275 90.860 46.445 90.880 ;
        RECT 45.655 90.445 45.885 90.860 ;
        RECT 46.245 90.445 46.475 90.860 ;
        RECT 45.655 90.275 46.475 90.445 ;
        RECT 45.655 89.860 45.885 90.275 ;
        RECT 46.245 89.860 46.475 90.275 ;
        RECT 45.685 89.840 45.855 89.860 ;
        RECT 46.275 89.840 46.445 89.860 ;
        RECT 46.730 89.655 46.900 91.065 ;
        RECT 47.185 90.860 47.355 90.880 ;
        RECT 47.775 90.860 47.945 91.455 ;
        RECT 48.085 91.065 48.545 91.295 ;
        RECT 47.155 89.860 47.385 90.860 ;
        RECT 47.745 89.860 47.975 90.860 ;
        RECT 45.085 89.425 45.545 89.655 ;
        RECT 46.585 89.425 47.045 89.655 ;
        RECT 45.230 87.720 45.400 89.425 ;
        RECT 45.610 88.465 45.930 88.725 ;
        RECT 45.085 87.490 45.545 87.720 ;
        RECT 44.775 87.330 44.945 87.350 ;
        RECT 44.155 86.680 44.385 87.330 ;
        RECT 44.745 86.680 44.975 87.330 ;
        RECT 44.185 86.660 44.355 86.680 ;
        RECT 43.585 86.290 44.045 86.520 ;
        RECT 44.775 86.085 44.945 86.680 ;
        RECT 45.230 86.565 45.400 87.490 ;
        RECT 45.685 87.330 45.855 88.465 ;
        RECT 46.730 87.720 46.900 89.425 ;
        RECT 47.185 88.725 47.355 89.860 ;
        RECT 47.775 89.840 47.945 89.860 ;
        RECT 48.230 89.655 48.400 91.065 ;
        RECT 48.640 90.635 48.900 90.955 ;
        RECT 49.275 90.860 49.445 91.455 ;
        RECT 49.585 91.065 50.045 91.295 ;
        RECT 51.085 91.065 51.545 91.295 ;
        RECT 48.655 89.860 48.885 90.635 ;
        RECT 49.245 89.860 49.475 90.860 ;
        RECT 48.085 89.425 48.545 89.655 ;
        RECT 48.230 88.725 48.400 89.425 ;
        RECT 47.110 88.465 47.430 88.725 ;
        RECT 48.155 88.465 48.475 88.725 ;
        RECT 46.585 87.490 47.045 87.720 ;
        RECT 46.275 87.330 46.445 87.350 ;
        RECT 45.655 86.680 45.885 87.330 ;
        RECT 46.245 86.680 46.475 87.330 ;
        RECT 45.685 86.660 45.855 86.680 ;
        RECT 45.185 86.520 45.445 86.565 ;
        RECT 45.085 86.290 45.545 86.520 ;
        RECT 45.185 86.245 45.445 86.290 ;
        RECT 46.275 86.085 46.445 86.680 ;
        RECT 46.730 86.565 46.900 87.490 ;
        RECT 47.185 87.330 47.355 88.465 ;
        RECT 48.230 87.720 48.400 88.465 ;
        RECT 48.085 87.490 48.545 87.720 ;
        RECT 47.775 87.330 47.945 87.350 ;
        RECT 47.155 86.680 47.385 87.330 ;
        RECT 47.745 86.680 47.975 87.330 ;
        RECT 47.185 86.660 47.355 86.680 ;
        RECT 46.685 86.520 46.945 86.565 ;
        RECT 46.585 86.290 47.045 86.520 ;
        RECT 46.685 86.245 46.945 86.290 ;
        RECT 47.775 86.085 47.945 86.680 ;
        RECT 48.230 86.520 48.400 87.490 ;
        RECT 48.685 87.330 48.855 89.860 ;
        RECT 49.275 89.840 49.445 89.860 ;
        RECT 49.730 89.655 49.900 91.065 ;
        RECT 50.185 90.860 50.355 90.880 ;
        RECT 50.775 90.860 50.945 90.880 ;
        RECT 50.155 90.445 50.385 90.860 ;
        RECT 50.745 90.445 50.975 90.860 ;
        RECT 50.155 90.275 50.975 90.445 ;
        RECT 50.155 89.860 50.385 90.275 ;
        RECT 50.745 89.860 50.975 90.275 ;
        RECT 50.185 89.840 50.355 89.860 ;
        RECT 50.775 89.840 50.945 89.860 ;
        RECT 51.230 89.655 51.400 91.065 ;
        RECT 51.685 90.860 51.855 90.880 ;
        RECT 52.275 90.860 52.445 91.455 ;
        RECT 52.585 91.065 53.045 91.295 ;
        RECT 51.655 89.860 51.885 90.860 ;
        RECT 52.245 89.860 52.475 90.860 ;
        RECT 49.585 89.425 50.045 89.655 ;
        RECT 51.085 89.425 51.545 89.655 ;
        RECT 49.730 87.720 49.900 89.425 ;
        RECT 50.110 88.465 50.430 88.725 ;
        RECT 49.585 87.490 50.045 87.720 ;
        RECT 49.275 87.330 49.445 87.350 ;
        RECT 48.655 86.680 48.885 87.330 ;
        RECT 49.245 86.680 49.475 87.330 ;
        RECT 48.685 86.660 48.855 86.680 ;
        RECT 48.085 86.290 48.545 86.520 ;
        RECT 49.275 86.085 49.445 86.680 ;
        RECT 49.730 86.565 49.900 87.490 ;
        RECT 50.185 87.330 50.355 88.465 ;
        RECT 51.230 87.720 51.400 89.425 ;
        RECT 51.685 88.725 51.855 89.860 ;
        RECT 52.275 89.840 52.445 89.860 ;
        RECT 52.730 89.655 52.900 91.065 ;
        RECT 53.140 90.635 53.400 90.955 ;
        RECT 53.775 90.860 53.945 91.455 ;
        RECT 54.085 91.065 54.545 91.295 ;
        RECT 55.585 91.065 56.045 91.295 ;
        RECT 53.155 89.860 53.385 90.635 ;
        RECT 53.745 89.860 53.975 90.860 ;
        RECT 52.585 89.425 53.045 89.655 ;
        RECT 52.730 88.725 52.900 89.425 ;
        RECT 51.610 88.465 51.930 88.725 ;
        RECT 52.655 88.465 52.975 88.725 ;
        RECT 51.085 87.490 51.545 87.720 ;
        RECT 50.775 87.330 50.945 87.350 ;
        RECT 50.155 86.680 50.385 87.330 ;
        RECT 50.745 86.680 50.975 87.330 ;
        RECT 50.185 86.660 50.355 86.680 ;
        RECT 49.685 86.520 49.945 86.565 ;
        RECT 49.585 86.290 50.045 86.520 ;
        RECT 49.685 86.245 49.945 86.290 ;
        RECT 50.775 86.085 50.945 86.680 ;
        RECT 51.230 86.565 51.400 87.490 ;
        RECT 51.685 87.330 51.855 88.465 ;
        RECT 52.730 87.720 52.900 88.465 ;
        RECT 52.585 87.490 53.045 87.720 ;
        RECT 52.275 87.330 52.445 87.350 ;
        RECT 51.655 86.680 51.885 87.330 ;
        RECT 52.245 86.680 52.475 87.330 ;
        RECT 51.685 86.660 51.855 86.680 ;
        RECT 51.185 86.520 51.445 86.565 ;
        RECT 51.085 86.290 51.545 86.520 ;
        RECT 51.185 86.245 51.445 86.290 ;
        RECT 52.275 86.085 52.445 86.680 ;
        RECT 52.730 86.520 52.900 87.490 ;
        RECT 53.185 87.330 53.355 89.860 ;
        RECT 53.775 89.840 53.945 89.860 ;
        RECT 54.230 89.655 54.400 91.065 ;
        RECT 54.685 90.860 54.855 90.880 ;
        RECT 55.275 90.860 55.445 90.880 ;
        RECT 54.655 90.445 54.885 90.860 ;
        RECT 55.245 90.445 55.475 90.860 ;
        RECT 54.655 90.275 55.475 90.445 ;
        RECT 54.655 89.860 54.885 90.275 ;
        RECT 55.245 89.860 55.475 90.275 ;
        RECT 54.685 89.840 54.855 89.860 ;
        RECT 55.275 89.840 55.445 89.860 ;
        RECT 55.730 89.655 55.900 91.065 ;
        RECT 56.185 90.860 56.355 90.880 ;
        RECT 56.775 90.860 56.945 91.455 ;
        RECT 57.085 91.065 57.545 91.295 ;
        RECT 56.155 89.860 56.385 90.860 ;
        RECT 56.745 89.860 56.975 90.860 ;
        RECT 54.085 89.425 54.545 89.655 ;
        RECT 55.585 89.425 56.045 89.655 ;
        RECT 54.230 87.720 54.400 89.425 ;
        RECT 54.610 88.465 54.930 88.725 ;
        RECT 54.085 87.490 54.545 87.720 ;
        RECT 53.775 87.330 53.945 87.350 ;
        RECT 53.155 86.680 53.385 87.330 ;
        RECT 53.745 86.680 53.975 87.330 ;
        RECT 53.185 86.660 53.355 86.680 ;
        RECT 52.585 86.290 53.045 86.520 ;
        RECT 53.775 86.085 53.945 86.680 ;
        RECT 54.230 86.565 54.400 87.490 ;
        RECT 54.685 87.330 54.855 88.465 ;
        RECT 55.730 87.720 55.900 89.425 ;
        RECT 56.185 88.725 56.355 89.860 ;
        RECT 56.775 89.840 56.945 89.860 ;
        RECT 57.230 89.655 57.400 91.065 ;
        RECT 57.640 90.635 57.900 90.955 ;
        RECT 58.275 90.860 58.445 91.455 ;
        RECT 58.585 91.065 59.045 91.295 ;
        RECT 60.085 91.065 60.545 91.295 ;
        RECT 57.655 89.860 57.885 90.635 ;
        RECT 58.245 89.860 58.475 90.860 ;
        RECT 57.085 89.425 57.545 89.655 ;
        RECT 57.230 88.725 57.400 89.425 ;
        RECT 56.110 88.465 56.430 88.725 ;
        RECT 57.155 88.465 57.475 88.725 ;
        RECT 55.585 87.490 56.045 87.720 ;
        RECT 55.275 87.330 55.445 87.350 ;
        RECT 54.655 86.680 54.885 87.330 ;
        RECT 55.245 86.680 55.475 87.330 ;
        RECT 54.685 86.660 54.855 86.680 ;
        RECT 54.185 86.520 54.445 86.565 ;
        RECT 54.085 86.290 54.545 86.520 ;
        RECT 54.185 86.245 54.445 86.290 ;
        RECT 55.275 86.085 55.445 86.680 ;
        RECT 55.730 86.565 55.900 87.490 ;
        RECT 56.185 87.330 56.355 88.465 ;
        RECT 57.230 87.720 57.400 88.465 ;
        RECT 57.085 87.490 57.545 87.720 ;
        RECT 56.775 87.330 56.945 87.350 ;
        RECT 56.155 86.680 56.385 87.330 ;
        RECT 56.745 86.680 56.975 87.330 ;
        RECT 56.185 86.660 56.355 86.680 ;
        RECT 55.685 86.520 55.945 86.565 ;
        RECT 55.585 86.290 56.045 86.520 ;
        RECT 55.685 86.245 55.945 86.290 ;
        RECT 56.775 86.085 56.945 86.680 ;
        RECT 57.230 86.520 57.400 87.490 ;
        RECT 57.685 87.330 57.855 89.860 ;
        RECT 58.275 89.840 58.445 89.860 ;
        RECT 58.730 89.655 58.900 91.065 ;
        RECT 59.185 90.860 59.355 90.880 ;
        RECT 59.775 90.860 59.945 90.880 ;
        RECT 59.155 90.445 59.385 90.860 ;
        RECT 59.745 90.445 59.975 90.860 ;
        RECT 59.155 90.275 59.975 90.445 ;
        RECT 59.155 89.860 59.385 90.275 ;
        RECT 59.745 89.860 59.975 90.275 ;
        RECT 59.185 89.840 59.355 89.860 ;
        RECT 59.775 89.840 59.945 89.860 ;
        RECT 60.230 89.655 60.400 91.065 ;
        RECT 60.685 90.860 60.855 90.880 ;
        RECT 61.275 90.860 61.445 91.455 ;
        RECT 61.585 91.065 62.045 91.295 ;
        RECT 60.655 89.860 60.885 90.860 ;
        RECT 61.245 89.860 61.475 90.860 ;
        RECT 58.585 89.425 59.045 89.655 ;
        RECT 60.085 89.425 60.545 89.655 ;
        RECT 58.730 87.720 58.900 89.425 ;
        RECT 59.110 88.465 59.430 88.725 ;
        RECT 58.585 87.490 59.045 87.720 ;
        RECT 58.275 87.330 58.445 87.350 ;
        RECT 57.655 86.680 57.885 87.330 ;
        RECT 58.245 86.680 58.475 87.330 ;
        RECT 57.685 86.660 57.855 86.680 ;
        RECT 57.085 86.290 57.545 86.520 ;
        RECT 58.275 86.085 58.445 86.680 ;
        RECT 58.730 86.565 58.900 87.490 ;
        RECT 59.185 87.330 59.355 88.465 ;
        RECT 60.230 87.720 60.400 89.425 ;
        RECT 60.685 88.725 60.855 89.860 ;
        RECT 61.275 89.840 61.445 89.860 ;
        RECT 61.730 89.655 61.900 91.065 ;
        RECT 62.140 90.635 62.400 90.955 ;
        RECT 62.775 90.860 62.945 91.455 ;
        RECT 63.085 91.065 63.545 91.295 ;
        RECT 64.585 91.065 65.045 91.295 ;
        RECT 62.155 89.860 62.385 90.635 ;
        RECT 62.745 89.860 62.975 90.860 ;
        RECT 61.585 89.425 62.045 89.655 ;
        RECT 61.730 88.725 61.900 89.425 ;
        RECT 60.610 88.465 60.930 88.725 ;
        RECT 61.655 88.465 61.975 88.725 ;
        RECT 60.085 87.490 60.545 87.720 ;
        RECT 59.775 87.330 59.945 87.350 ;
        RECT 59.155 86.680 59.385 87.330 ;
        RECT 59.745 86.680 59.975 87.330 ;
        RECT 59.185 86.660 59.355 86.680 ;
        RECT 58.685 86.520 58.945 86.565 ;
        RECT 58.585 86.290 59.045 86.520 ;
        RECT 58.685 86.245 58.945 86.290 ;
        RECT 59.775 86.085 59.945 86.680 ;
        RECT 60.230 86.565 60.400 87.490 ;
        RECT 60.685 87.330 60.855 88.465 ;
        RECT 61.730 87.720 61.900 88.465 ;
        RECT 61.585 87.490 62.045 87.720 ;
        RECT 61.275 87.330 61.445 87.350 ;
        RECT 60.655 86.680 60.885 87.330 ;
        RECT 61.245 86.680 61.475 87.330 ;
        RECT 60.685 86.660 60.855 86.680 ;
        RECT 60.185 86.520 60.445 86.565 ;
        RECT 60.085 86.290 60.545 86.520 ;
        RECT 60.185 86.245 60.445 86.290 ;
        RECT 61.275 86.085 61.445 86.680 ;
        RECT 61.730 86.520 61.900 87.490 ;
        RECT 62.185 87.330 62.355 89.860 ;
        RECT 62.775 89.840 62.945 89.860 ;
        RECT 63.230 89.655 63.400 91.065 ;
        RECT 63.685 90.860 63.855 90.880 ;
        RECT 64.275 90.860 64.445 90.880 ;
        RECT 63.655 90.445 63.885 90.860 ;
        RECT 64.245 90.445 64.475 90.860 ;
        RECT 63.655 90.275 64.475 90.445 ;
        RECT 63.655 89.860 63.885 90.275 ;
        RECT 64.245 89.860 64.475 90.275 ;
        RECT 63.685 89.840 63.855 89.860 ;
        RECT 64.275 89.840 64.445 89.860 ;
        RECT 64.730 89.655 64.900 91.065 ;
        RECT 65.185 90.860 65.355 90.880 ;
        RECT 65.775 90.860 65.945 91.455 ;
        RECT 66.085 91.065 66.545 91.295 ;
        RECT 65.155 89.860 65.385 90.860 ;
        RECT 65.745 89.860 65.975 90.860 ;
        RECT 63.085 89.425 63.545 89.655 ;
        RECT 64.585 89.425 65.045 89.655 ;
        RECT 63.230 87.720 63.400 89.425 ;
        RECT 63.610 88.465 63.930 88.725 ;
        RECT 63.085 87.490 63.545 87.720 ;
        RECT 62.775 87.330 62.945 87.350 ;
        RECT 62.155 86.680 62.385 87.330 ;
        RECT 62.745 86.680 62.975 87.330 ;
        RECT 62.185 86.660 62.355 86.680 ;
        RECT 61.585 86.290 62.045 86.520 ;
        RECT 62.775 86.085 62.945 86.680 ;
        RECT 63.230 86.565 63.400 87.490 ;
        RECT 63.685 87.330 63.855 88.465 ;
        RECT 64.730 87.720 64.900 89.425 ;
        RECT 65.185 88.725 65.355 89.860 ;
        RECT 65.775 89.840 65.945 89.860 ;
        RECT 66.230 89.655 66.400 91.065 ;
        RECT 66.640 90.635 66.900 90.955 ;
        RECT 67.275 90.860 67.445 91.455 ;
        RECT 67.585 91.065 68.045 91.295 ;
        RECT 69.085 91.065 69.545 91.295 ;
        RECT 66.655 89.860 66.885 90.635 ;
        RECT 67.245 89.860 67.475 90.860 ;
        RECT 66.085 89.425 66.545 89.655 ;
        RECT 66.230 88.725 66.400 89.425 ;
        RECT 65.110 88.465 65.430 88.725 ;
        RECT 66.155 88.465 66.475 88.725 ;
        RECT 64.585 87.490 65.045 87.720 ;
        RECT 64.275 87.330 64.445 87.350 ;
        RECT 63.655 86.680 63.885 87.330 ;
        RECT 64.245 86.680 64.475 87.330 ;
        RECT 63.685 86.660 63.855 86.680 ;
        RECT 63.185 86.520 63.445 86.565 ;
        RECT 63.085 86.290 63.545 86.520 ;
        RECT 63.185 86.245 63.445 86.290 ;
        RECT 64.275 86.085 64.445 86.680 ;
        RECT 64.730 86.565 64.900 87.490 ;
        RECT 65.185 87.330 65.355 88.465 ;
        RECT 66.230 87.720 66.400 88.465 ;
        RECT 66.085 87.490 66.545 87.720 ;
        RECT 65.775 87.330 65.945 87.350 ;
        RECT 65.155 86.680 65.385 87.330 ;
        RECT 65.745 86.680 65.975 87.330 ;
        RECT 65.185 86.660 65.355 86.680 ;
        RECT 64.685 86.520 64.945 86.565 ;
        RECT 64.585 86.290 65.045 86.520 ;
        RECT 64.685 86.245 64.945 86.290 ;
        RECT 65.775 86.085 65.945 86.680 ;
        RECT 66.230 86.520 66.400 87.490 ;
        RECT 66.685 87.330 66.855 89.860 ;
        RECT 67.275 89.840 67.445 89.860 ;
        RECT 67.730 89.655 67.900 91.065 ;
        RECT 68.185 90.860 68.355 90.880 ;
        RECT 68.775 90.860 68.945 90.880 ;
        RECT 68.155 90.445 68.385 90.860 ;
        RECT 68.745 90.445 68.975 90.860 ;
        RECT 68.155 90.275 68.975 90.445 ;
        RECT 68.155 89.860 68.385 90.275 ;
        RECT 68.745 89.860 68.975 90.275 ;
        RECT 68.185 89.840 68.355 89.860 ;
        RECT 68.775 89.840 68.945 89.860 ;
        RECT 69.230 89.655 69.400 91.065 ;
        RECT 69.685 90.860 69.855 90.880 ;
        RECT 70.275 90.860 70.445 91.455 ;
        RECT 70.585 91.065 71.045 91.295 ;
        RECT 69.655 89.860 69.885 90.860 ;
        RECT 70.245 89.860 70.475 90.860 ;
        RECT 67.585 89.425 68.045 89.655 ;
        RECT 69.085 89.425 69.545 89.655 ;
        RECT 67.730 87.720 67.900 89.425 ;
        RECT 68.110 88.465 68.430 88.725 ;
        RECT 67.585 87.490 68.045 87.720 ;
        RECT 67.275 87.330 67.445 87.350 ;
        RECT 66.655 86.680 66.885 87.330 ;
        RECT 67.245 86.680 67.475 87.330 ;
        RECT 66.685 86.660 66.855 86.680 ;
        RECT 66.085 86.290 66.545 86.520 ;
        RECT 67.275 86.085 67.445 86.680 ;
        RECT 67.730 86.565 67.900 87.490 ;
        RECT 68.185 87.330 68.355 88.465 ;
        RECT 69.230 87.720 69.400 89.425 ;
        RECT 69.685 88.725 69.855 89.860 ;
        RECT 70.275 89.840 70.445 89.860 ;
        RECT 70.730 89.655 70.900 91.065 ;
        RECT 71.140 90.635 71.400 90.955 ;
        RECT 71.775 90.860 71.945 91.455 ;
        RECT 72.085 91.065 72.545 91.295 ;
        RECT 73.585 91.065 74.045 91.295 ;
        RECT 71.155 89.860 71.385 90.635 ;
        RECT 71.745 89.860 71.975 90.860 ;
        RECT 70.585 89.425 71.045 89.655 ;
        RECT 70.730 88.725 70.900 89.425 ;
        RECT 69.610 88.465 69.930 88.725 ;
        RECT 70.655 88.465 70.975 88.725 ;
        RECT 69.085 87.490 69.545 87.720 ;
        RECT 68.775 87.330 68.945 87.350 ;
        RECT 68.155 86.680 68.385 87.330 ;
        RECT 68.745 86.680 68.975 87.330 ;
        RECT 68.185 86.660 68.355 86.680 ;
        RECT 67.685 86.520 67.945 86.565 ;
        RECT 67.585 86.290 68.045 86.520 ;
        RECT 67.685 86.245 67.945 86.290 ;
        RECT 68.775 86.085 68.945 86.680 ;
        RECT 69.230 86.565 69.400 87.490 ;
        RECT 69.685 87.330 69.855 88.465 ;
        RECT 70.730 87.720 70.900 88.465 ;
        RECT 70.585 87.490 71.045 87.720 ;
        RECT 70.275 87.330 70.445 87.350 ;
        RECT 69.655 86.680 69.885 87.330 ;
        RECT 70.245 86.680 70.475 87.330 ;
        RECT 69.685 86.660 69.855 86.680 ;
        RECT 69.185 86.520 69.445 86.565 ;
        RECT 69.085 86.290 69.545 86.520 ;
        RECT 69.185 86.245 69.445 86.290 ;
        RECT 70.275 86.085 70.445 86.680 ;
        RECT 70.730 86.520 70.900 87.490 ;
        RECT 71.185 87.330 71.355 89.860 ;
        RECT 71.775 89.840 71.945 89.860 ;
        RECT 72.230 89.655 72.400 91.065 ;
        RECT 72.685 90.860 72.855 90.880 ;
        RECT 73.275 90.860 73.445 90.880 ;
        RECT 72.655 90.445 72.885 90.860 ;
        RECT 73.245 90.445 73.475 90.860 ;
        RECT 72.655 90.275 73.475 90.445 ;
        RECT 72.655 89.860 72.885 90.275 ;
        RECT 73.245 89.860 73.475 90.275 ;
        RECT 72.685 89.840 72.855 89.860 ;
        RECT 73.275 89.840 73.445 89.860 ;
        RECT 73.730 89.655 73.900 91.065 ;
        RECT 74.185 90.860 74.355 90.880 ;
        RECT 74.775 90.860 74.945 91.455 ;
        RECT 75.085 91.065 75.545 91.295 ;
        RECT 74.155 89.860 74.385 90.860 ;
        RECT 74.745 89.860 74.975 90.860 ;
        RECT 72.085 89.425 72.545 89.655 ;
        RECT 73.585 89.425 74.045 89.655 ;
        RECT 72.230 87.720 72.400 89.425 ;
        RECT 72.610 88.465 72.930 88.725 ;
        RECT 72.085 87.490 72.545 87.720 ;
        RECT 71.775 87.330 71.945 87.350 ;
        RECT 71.155 86.680 71.385 87.330 ;
        RECT 71.745 86.680 71.975 87.330 ;
        RECT 71.185 86.660 71.355 86.680 ;
        RECT 70.585 86.290 71.045 86.520 ;
        RECT 71.775 86.085 71.945 86.680 ;
        RECT 72.230 86.565 72.400 87.490 ;
        RECT 72.685 87.330 72.855 88.465 ;
        RECT 73.730 87.720 73.900 89.425 ;
        RECT 74.185 88.725 74.355 89.860 ;
        RECT 74.775 89.840 74.945 89.860 ;
        RECT 75.230 89.655 75.400 91.065 ;
        RECT 75.640 90.635 75.900 90.955 ;
        RECT 76.275 90.860 76.445 91.455 ;
        RECT 76.585 91.065 77.045 91.295 ;
        RECT 78.085 91.065 78.545 91.295 ;
        RECT 75.655 89.860 75.885 90.635 ;
        RECT 76.245 89.860 76.475 90.860 ;
        RECT 75.085 89.425 75.545 89.655 ;
        RECT 75.230 88.725 75.400 89.425 ;
        RECT 74.110 88.465 74.430 88.725 ;
        RECT 75.155 88.465 75.475 88.725 ;
        RECT 73.585 87.490 74.045 87.720 ;
        RECT 73.275 87.330 73.445 87.350 ;
        RECT 72.655 86.680 72.885 87.330 ;
        RECT 73.245 86.680 73.475 87.330 ;
        RECT 72.685 86.660 72.855 86.680 ;
        RECT 72.185 86.520 72.445 86.565 ;
        RECT 72.085 86.290 72.545 86.520 ;
        RECT 72.185 86.245 72.445 86.290 ;
        RECT 73.275 86.085 73.445 86.680 ;
        RECT 73.730 86.565 73.900 87.490 ;
        RECT 74.185 87.330 74.355 88.465 ;
        RECT 75.230 87.720 75.400 88.465 ;
        RECT 75.085 87.490 75.545 87.720 ;
        RECT 74.775 87.330 74.945 87.350 ;
        RECT 74.155 86.680 74.385 87.330 ;
        RECT 74.745 86.680 74.975 87.330 ;
        RECT 74.185 86.660 74.355 86.680 ;
        RECT 73.685 86.520 73.945 86.565 ;
        RECT 73.585 86.290 74.045 86.520 ;
        RECT 73.685 86.245 73.945 86.290 ;
        RECT 74.775 86.085 74.945 86.680 ;
        RECT 75.230 86.520 75.400 87.490 ;
        RECT 75.685 87.330 75.855 89.860 ;
        RECT 76.275 89.840 76.445 89.860 ;
        RECT 76.730 89.655 76.900 91.065 ;
        RECT 77.185 90.860 77.355 90.880 ;
        RECT 77.775 90.860 77.945 90.880 ;
        RECT 77.155 90.445 77.385 90.860 ;
        RECT 77.745 90.445 77.975 90.860 ;
        RECT 77.155 90.275 77.975 90.445 ;
        RECT 77.155 89.860 77.385 90.275 ;
        RECT 77.745 89.860 77.975 90.275 ;
        RECT 77.185 89.840 77.355 89.860 ;
        RECT 77.775 89.840 77.945 89.860 ;
        RECT 78.230 89.655 78.400 91.065 ;
        RECT 78.685 90.860 78.855 90.880 ;
        RECT 79.275 90.860 79.445 91.455 ;
        RECT 79.585 91.065 80.045 91.295 ;
        RECT 78.655 89.860 78.885 90.860 ;
        RECT 79.245 89.860 79.475 90.860 ;
        RECT 76.585 89.425 77.045 89.655 ;
        RECT 78.085 89.425 78.545 89.655 ;
        RECT 76.730 87.720 76.900 89.425 ;
        RECT 77.110 88.465 77.430 88.725 ;
        RECT 76.585 87.490 77.045 87.720 ;
        RECT 76.275 87.330 76.445 87.350 ;
        RECT 75.655 86.680 75.885 87.330 ;
        RECT 76.245 86.680 76.475 87.330 ;
        RECT 75.685 86.660 75.855 86.680 ;
        RECT 75.085 86.290 75.545 86.520 ;
        RECT 76.275 86.085 76.445 86.680 ;
        RECT 76.730 86.565 76.900 87.490 ;
        RECT 77.185 87.330 77.355 88.465 ;
        RECT 78.230 87.720 78.400 89.425 ;
        RECT 78.685 88.725 78.855 89.860 ;
        RECT 79.275 89.840 79.445 89.860 ;
        RECT 79.730 89.655 79.900 91.065 ;
        RECT 80.140 90.635 80.400 90.955 ;
        RECT 80.775 90.860 80.945 91.455 ;
        RECT 81.085 91.065 81.545 91.295 ;
        RECT 82.585 91.065 83.045 91.295 ;
        RECT 80.155 89.860 80.385 90.635 ;
        RECT 80.745 89.860 80.975 90.860 ;
        RECT 79.585 89.425 80.045 89.655 ;
        RECT 79.730 88.725 79.900 89.425 ;
        RECT 78.610 88.465 78.930 88.725 ;
        RECT 79.655 88.465 79.975 88.725 ;
        RECT 78.085 87.490 78.545 87.720 ;
        RECT 77.775 87.330 77.945 87.350 ;
        RECT 77.155 86.680 77.385 87.330 ;
        RECT 77.745 86.680 77.975 87.330 ;
        RECT 77.185 86.660 77.355 86.680 ;
        RECT 76.685 86.520 76.945 86.565 ;
        RECT 76.585 86.290 77.045 86.520 ;
        RECT 76.685 86.245 76.945 86.290 ;
        RECT 77.775 86.085 77.945 86.680 ;
        RECT 78.230 86.565 78.400 87.490 ;
        RECT 78.685 87.330 78.855 88.465 ;
        RECT 79.730 87.720 79.900 88.465 ;
        RECT 79.585 87.490 80.045 87.720 ;
        RECT 79.275 87.330 79.445 87.350 ;
        RECT 78.655 86.680 78.885 87.330 ;
        RECT 79.245 86.680 79.475 87.330 ;
        RECT 78.685 86.660 78.855 86.680 ;
        RECT 78.185 86.520 78.445 86.565 ;
        RECT 78.085 86.290 78.545 86.520 ;
        RECT 78.185 86.245 78.445 86.290 ;
        RECT 79.275 86.085 79.445 86.680 ;
        RECT 79.730 86.520 79.900 87.490 ;
        RECT 80.185 87.330 80.355 89.860 ;
        RECT 80.775 89.840 80.945 89.860 ;
        RECT 81.230 89.655 81.400 91.065 ;
        RECT 81.685 90.860 81.855 90.880 ;
        RECT 82.275 90.860 82.445 90.880 ;
        RECT 81.655 90.445 81.885 90.860 ;
        RECT 82.245 90.445 82.475 90.860 ;
        RECT 81.655 90.275 82.475 90.445 ;
        RECT 81.655 89.860 81.885 90.275 ;
        RECT 82.245 89.860 82.475 90.275 ;
        RECT 81.685 89.840 81.855 89.860 ;
        RECT 82.275 89.840 82.445 89.860 ;
        RECT 82.730 89.655 82.900 91.065 ;
        RECT 83.185 90.860 83.355 90.880 ;
        RECT 83.775 90.860 83.945 91.455 ;
        RECT 84.085 91.065 84.545 91.295 ;
        RECT 83.155 89.860 83.385 90.860 ;
        RECT 83.745 89.860 83.975 90.860 ;
        RECT 81.085 89.425 81.545 89.655 ;
        RECT 82.585 89.425 83.045 89.655 ;
        RECT 81.230 87.720 81.400 89.425 ;
        RECT 81.610 88.465 81.930 88.725 ;
        RECT 81.085 87.490 81.545 87.720 ;
        RECT 80.775 87.330 80.945 87.350 ;
        RECT 80.155 86.680 80.385 87.330 ;
        RECT 80.745 86.680 80.975 87.330 ;
        RECT 80.185 86.660 80.355 86.680 ;
        RECT 79.585 86.290 80.045 86.520 ;
        RECT 80.775 86.085 80.945 86.680 ;
        RECT 81.230 86.565 81.400 87.490 ;
        RECT 81.685 87.330 81.855 88.465 ;
        RECT 82.730 87.720 82.900 89.425 ;
        RECT 83.185 88.725 83.355 89.860 ;
        RECT 83.775 89.840 83.945 89.860 ;
        RECT 84.230 89.655 84.400 91.065 ;
        RECT 84.640 90.635 84.900 90.955 ;
        RECT 85.275 90.860 85.445 91.455 ;
        RECT 85.585 91.065 86.045 91.295 ;
        RECT 87.085 91.065 87.545 91.295 ;
        RECT 84.655 89.860 84.885 90.635 ;
        RECT 85.245 89.860 85.475 90.860 ;
        RECT 84.085 89.425 84.545 89.655 ;
        RECT 84.230 88.725 84.400 89.425 ;
        RECT 83.110 88.465 83.430 88.725 ;
        RECT 84.155 88.465 84.475 88.725 ;
        RECT 82.585 87.490 83.045 87.720 ;
        RECT 82.275 87.330 82.445 87.350 ;
        RECT 81.655 86.680 81.885 87.330 ;
        RECT 82.245 86.680 82.475 87.330 ;
        RECT 81.685 86.660 81.855 86.680 ;
        RECT 81.185 86.520 81.445 86.565 ;
        RECT 81.085 86.290 81.545 86.520 ;
        RECT 81.185 86.245 81.445 86.290 ;
        RECT 82.275 86.085 82.445 86.680 ;
        RECT 82.730 86.565 82.900 87.490 ;
        RECT 83.185 87.330 83.355 88.465 ;
        RECT 84.230 87.720 84.400 88.465 ;
        RECT 84.085 87.490 84.545 87.720 ;
        RECT 83.775 87.330 83.945 87.350 ;
        RECT 83.155 86.680 83.385 87.330 ;
        RECT 83.745 86.680 83.975 87.330 ;
        RECT 83.185 86.660 83.355 86.680 ;
        RECT 82.685 86.520 82.945 86.565 ;
        RECT 82.585 86.290 83.045 86.520 ;
        RECT 82.685 86.245 82.945 86.290 ;
        RECT 83.775 86.085 83.945 86.680 ;
        RECT 84.230 86.520 84.400 87.490 ;
        RECT 84.685 87.330 84.855 89.860 ;
        RECT 85.275 89.840 85.445 89.860 ;
        RECT 85.730 89.655 85.900 91.065 ;
        RECT 86.185 90.860 86.355 90.880 ;
        RECT 86.775 90.860 86.945 90.880 ;
        RECT 86.155 90.445 86.385 90.860 ;
        RECT 86.745 90.445 86.975 90.860 ;
        RECT 86.155 90.275 86.975 90.445 ;
        RECT 86.155 89.860 86.385 90.275 ;
        RECT 86.745 89.860 86.975 90.275 ;
        RECT 86.185 89.840 86.355 89.860 ;
        RECT 86.775 89.840 86.945 89.860 ;
        RECT 87.230 89.655 87.400 91.065 ;
        RECT 87.685 90.860 87.855 90.880 ;
        RECT 88.275 90.860 88.445 91.455 ;
        RECT 88.585 91.065 89.045 91.295 ;
        RECT 87.655 89.860 87.885 90.860 ;
        RECT 88.245 89.860 88.475 90.860 ;
        RECT 85.585 89.425 86.045 89.655 ;
        RECT 87.085 89.425 87.545 89.655 ;
        RECT 85.730 87.720 85.900 89.425 ;
        RECT 86.110 88.465 86.430 88.725 ;
        RECT 85.585 87.490 86.045 87.720 ;
        RECT 85.275 87.330 85.445 87.350 ;
        RECT 84.655 86.680 84.885 87.330 ;
        RECT 85.245 86.680 85.475 87.330 ;
        RECT 84.685 86.660 84.855 86.680 ;
        RECT 84.085 86.290 84.545 86.520 ;
        RECT 85.275 86.085 85.445 86.680 ;
        RECT 85.730 86.565 85.900 87.490 ;
        RECT 86.185 87.330 86.355 88.465 ;
        RECT 87.230 87.720 87.400 89.425 ;
        RECT 87.685 88.725 87.855 89.860 ;
        RECT 88.275 89.840 88.445 89.860 ;
        RECT 88.730 89.655 88.900 91.065 ;
        RECT 89.140 90.635 89.400 90.955 ;
        RECT 89.775 90.860 89.945 91.455 ;
        RECT 90.085 91.065 90.545 91.295 ;
        RECT 91.585 91.065 92.045 91.295 ;
        RECT 89.155 89.860 89.385 90.635 ;
        RECT 89.745 89.860 89.975 90.860 ;
        RECT 88.585 89.425 89.045 89.655 ;
        RECT 88.730 88.725 88.900 89.425 ;
        RECT 87.610 88.465 87.930 88.725 ;
        RECT 88.655 88.465 88.975 88.725 ;
        RECT 87.085 87.490 87.545 87.720 ;
        RECT 86.775 87.330 86.945 87.350 ;
        RECT 86.155 86.680 86.385 87.330 ;
        RECT 86.745 86.680 86.975 87.330 ;
        RECT 86.185 86.660 86.355 86.680 ;
        RECT 85.685 86.520 85.945 86.565 ;
        RECT 85.585 86.290 86.045 86.520 ;
        RECT 85.685 86.245 85.945 86.290 ;
        RECT 86.775 86.085 86.945 86.680 ;
        RECT 87.230 86.565 87.400 87.490 ;
        RECT 87.685 87.330 87.855 88.465 ;
        RECT 88.730 87.720 88.900 88.465 ;
        RECT 88.585 87.490 89.045 87.720 ;
        RECT 88.275 87.330 88.445 87.350 ;
        RECT 87.655 86.680 87.885 87.330 ;
        RECT 88.245 86.680 88.475 87.330 ;
        RECT 87.685 86.660 87.855 86.680 ;
        RECT 87.185 86.520 87.445 86.565 ;
        RECT 87.085 86.290 87.545 86.520 ;
        RECT 87.185 86.245 87.445 86.290 ;
        RECT 88.275 86.085 88.445 86.680 ;
        RECT 88.730 86.520 88.900 87.490 ;
        RECT 89.185 87.330 89.355 89.860 ;
        RECT 89.775 89.840 89.945 89.860 ;
        RECT 90.230 89.655 90.400 91.065 ;
        RECT 90.685 90.860 90.855 90.880 ;
        RECT 91.275 90.860 91.445 90.880 ;
        RECT 90.655 90.445 90.885 90.860 ;
        RECT 91.245 90.445 91.475 90.860 ;
        RECT 90.655 90.275 91.475 90.445 ;
        RECT 90.655 89.860 90.885 90.275 ;
        RECT 91.245 89.860 91.475 90.275 ;
        RECT 90.685 89.840 90.855 89.860 ;
        RECT 91.275 89.840 91.445 89.860 ;
        RECT 91.730 89.655 91.900 91.065 ;
        RECT 92.185 90.860 92.355 90.880 ;
        RECT 92.775 90.860 92.945 91.455 ;
        RECT 93.085 91.065 93.545 91.295 ;
        RECT 92.155 89.860 92.385 90.860 ;
        RECT 92.745 89.860 92.975 90.860 ;
        RECT 90.085 89.425 90.545 89.655 ;
        RECT 91.585 89.425 92.045 89.655 ;
        RECT 90.230 87.720 90.400 89.425 ;
        RECT 90.610 88.465 90.930 88.725 ;
        RECT 90.085 87.490 90.545 87.720 ;
        RECT 89.775 87.330 89.945 87.350 ;
        RECT 89.155 86.680 89.385 87.330 ;
        RECT 89.745 86.680 89.975 87.330 ;
        RECT 89.185 86.660 89.355 86.680 ;
        RECT 88.585 86.290 89.045 86.520 ;
        RECT 89.775 86.085 89.945 86.680 ;
        RECT 90.230 86.565 90.400 87.490 ;
        RECT 90.685 87.330 90.855 88.465 ;
        RECT 91.730 87.720 91.900 89.425 ;
        RECT 92.185 88.725 92.355 89.860 ;
        RECT 92.775 89.840 92.945 89.860 ;
        RECT 93.230 89.655 93.400 91.065 ;
        RECT 93.640 90.635 93.900 90.955 ;
        RECT 94.275 90.860 94.445 91.455 ;
        RECT 94.585 91.065 95.045 91.295 ;
        RECT 96.085 91.065 96.545 91.295 ;
        RECT 93.655 89.860 93.885 90.635 ;
        RECT 94.245 89.860 94.475 90.860 ;
        RECT 93.085 89.425 93.545 89.655 ;
        RECT 93.230 88.725 93.400 89.425 ;
        RECT 92.110 88.465 92.430 88.725 ;
        RECT 93.155 88.465 93.475 88.725 ;
        RECT 91.585 87.490 92.045 87.720 ;
        RECT 91.275 87.330 91.445 87.350 ;
        RECT 90.655 86.680 90.885 87.330 ;
        RECT 91.245 86.680 91.475 87.330 ;
        RECT 90.685 86.660 90.855 86.680 ;
        RECT 90.185 86.520 90.445 86.565 ;
        RECT 90.085 86.290 90.545 86.520 ;
        RECT 90.185 86.245 90.445 86.290 ;
        RECT 91.275 86.085 91.445 86.680 ;
        RECT 91.730 86.565 91.900 87.490 ;
        RECT 92.185 87.330 92.355 88.465 ;
        RECT 93.230 87.720 93.400 88.465 ;
        RECT 93.085 87.490 93.545 87.720 ;
        RECT 92.775 87.330 92.945 87.350 ;
        RECT 92.155 86.680 92.385 87.330 ;
        RECT 92.745 86.680 92.975 87.330 ;
        RECT 92.185 86.660 92.355 86.680 ;
        RECT 91.685 86.520 91.945 86.565 ;
        RECT 91.585 86.290 92.045 86.520 ;
        RECT 91.685 86.245 91.945 86.290 ;
        RECT 92.775 86.085 92.945 86.680 ;
        RECT 93.230 86.520 93.400 87.490 ;
        RECT 93.685 87.330 93.855 89.860 ;
        RECT 94.275 89.840 94.445 89.860 ;
        RECT 94.730 89.655 94.900 91.065 ;
        RECT 95.185 90.860 95.355 90.880 ;
        RECT 95.775 90.860 95.945 90.880 ;
        RECT 95.155 90.445 95.385 90.860 ;
        RECT 95.745 90.445 95.975 90.860 ;
        RECT 95.155 90.275 95.975 90.445 ;
        RECT 95.155 89.860 95.385 90.275 ;
        RECT 95.745 89.860 95.975 90.275 ;
        RECT 95.185 89.840 95.355 89.860 ;
        RECT 95.775 89.840 95.945 89.860 ;
        RECT 96.230 89.655 96.400 91.065 ;
        RECT 96.685 90.860 96.855 90.880 ;
        RECT 97.275 90.860 97.445 91.455 ;
        RECT 97.585 91.065 98.045 91.295 ;
        RECT 96.655 89.860 96.885 90.860 ;
        RECT 97.245 89.860 97.475 90.860 ;
        RECT 94.585 89.425 95.045 89.655 ;
        RECT 96.085 89.425 96.545 89.655 ;
        RECT 94.730 87.720 94.900 89.425 ;
        RECT 95.110 88.465 95.430 88.725 ;
        RECT 94.585 87.490 95.045 87.720 ;
        RECT 94.275 87.330 94.445 87.350 ;
        RECT 93.655 86.680 93.885 87.330 ;
        RECT 94.245 86.680 94.475 87.330 ;
        RECT 93.685 86.660 93.855 86.680 ;
        RECT 93.085 86.290 93.545 86.520 ;
        RECT 94.275 86.085 94.445 86.680 ;
        RECT 94.730 86.565 94.900 87.490 ;
        RECT 95.185 87.330 95.355 88.465 ;
        RECT 96.230 87.720 96.400 89.425 ;
        RECT 96.685 88.725 96.855 89.860 ;
        RECT 97.275 89.840 97.445 89.860 ;
        RECT 97.730 89.655 97.900 91.065 ;
        RECT 98.140 90.635 98.400 90.955 ;
        RECT 98.775 90.860 98.945 91.455 ;
        RECT 99.085 91.065 99.545 91.295 ;
        RECT 100.585 91.065 101.045 91.295 ;
        RECT 98.155 89.860 98.385 90.635 ;
        RECT 98.745 89.860 98.975 90.860 ;
        RECT 97.585 89.425 98.045 89.655 ;
        RECT 97.730 88.725 97.900 89.425 ;
        RECT 96.610 88.465 96.930 88.725 ;
        RECT 97.655 88.465 97.975 88.725 ;
        RECT 96.085 87.490 96.545 87.720 ;
        RECT 95.775 87.330 95.945 87.350 ;
        RECT 95.155 86.680 95.385 87.330 ;
        RECT 95.745 86.680 95.975 87.330 ;
        RECT 95.185 86.660 95.355 86.680 ;
        RECT 94.685 86.520 94.945 86.565 ;
        RECT 94.585 86.290 95.045 86.520 ;
        RECT 94.685 86.245 94.945 86.290 ;
        RECT 95.775 86.085 95.945 86.680 ;
        RECT 96.230 86.565 96.400 87.490 ;
        RECT 96.685 87.330 96.855 88.465 ;
        RECT 97.730 87.720 97.900 88.465 ;
        RECT 97.585 87.490 98.045 87.720 ;
        RECT 97.275 87.330 97.445 87.350 ;
        RECT 96.655 86.680 96.885 87.330 ;
        RECT 97.245 86.680 97.475 87.330 ;
        RECT 96.685 86.660 96.855 86.680 ;
        RECT 96.185 86.520 96.445 86.565 ;
        RECT 96.085 86.290 96.545 86.520 ;
        RECT 96.185 86.245 96.445 86.290 ;
        RECT 97.275 86.085 97.445 86.680 ;
        RECT 97.730 86.520 97.900 87.490 ;
        RECT 98.185 87.330 98.355 89.860 ;
        RECT 98.775 89.840 98.945 89.860 ;
        RECT 99.230 89.655 99.400 91.065 ;
        RECT 99.685 90.860 99.855 90.880 ;
        RECT 100.275 90.860 100.445 90.880 ;
        RECT 99.655 90.445 99.885 90.860 ;
        RECT 100.245 90.445 100.475 90.860 ;
        RECT 99.655 90.275 100.475 90.445 ;
        RECT 99.655 89.860 99.885 90.275 ;
        RECT 100.245 89.860 100.475 90.275 ;
        RECT 99.685 89.840 99.855 89.860 ;
        RECT 100.275 89.840 100.445 89.860 ;
        RECT 100.730 89.655 100.900 91.065 ;
        RECT 101.185 90.860 101.355 90.880 ;
        RECT 101.775 90.860 101.945 91.455 ;
        RECT 102.085 91.065 102.545 91.295 ;
        RECT 101.155 89.860 101.385 90.860 ;
        RECT 101.745 89.860 101.975 90.860 ;
        RECT 99.085 89.425 99.545 89.655 ;
        RECT 100.585 89.425 101.045 89.655 ;
        RECT 99.230 87.720 99.400 89.425 ;
        RECT 99.610 88.465 99.930 88.725 ;
        RECT 99.085 87.490 99.545 87.720 ;
        RECT 98.775 87.330 98.945 87.350 ;
        RECT 98.155 86.680 98.385 87.330 ;
        RECT 98.745 86.680 98.975 87.330 ;
        RECT 98.185 86.660 98.355 86.680 ;
        RECT 97.585 86.290 98.045 86.520 ;
        RECT 98.775 86.085 98.945 86.680 ;
        RECT 99.230 86.565 99.400 87.490 ;
        RECT 99.685 87.330 99.855 88.465 ;
        RECT 100.730 87.720 100.900 89.425 ;
        RECT 101.185 88.725 101.355 89.860 ;
        RECT 101.775 89.840 101.945 89.860 ;
        RECT 102.230 89.655 102.400 91.065 ;
        RECT 102.640 90.635 102.900 90.955 ;
        RECT 103.275 90.860 103.445 91.455 ;
        RECT 103.585 91.065 104.045 91.295 ;
        RECT 105.085 91.065 105.545 91.295 ;
        RECT 102.655 89.860 102.885 90.635 ;
        RECT 103.245 89.860 103.475 90.860 ;
        RECT 102.085 89.425 102.545 89.655 ;
        RECT 102.230 88.725 102.400 89.425 ;
        RECT 101.110 88.465 101.430 88.725 ;
        RECT 102.155 88.465 102.475 88.725 ;
        RECT 100.585 87.490 101.045 87.720 ;
        RECT 100.275 87.330 100.445 87.350 ;
        RECT 99.655 86.680 99.885 87.330 ;
        RECT 100.245 86.680 100.475 87.330 ;
        RECT 99.685 86.660 99.855 86.680 ;
        RECT 99.185 86.520 99.445 86.565 ;
        RECT 99.085 86.290 99.545 86.520 ;
        RECT 99.185 86.245 99.445 86.290 ;
        RECT 100.275 86.085 100.445 86.680 ;
        RECT 100.730 86.565 100.900 87.490 ;
        RECT 101.185 87.330 101.355 88.465 ;
        RECT 102.230 87.720 102.400 88.465 ;
        RECT 102.085 87.490 102.545 87.720 ;
        RECT 101.775 87.330 101.945 87.350 ;
        RECT 101.155 86.680 101.385 87.330 ;
        RECT 101.745 86.680 101.975 87.330 ;
        RECT 101.185 86.660 101.355 86.680 ;
        RECT 100.685 86.520 100.945 86.565 ;
        RECT 100.585 86.290 101.045 86.520 ;
        RECT 100.685 86.245 100.945 86.290 ;
        RECT 101.775 86.085 101.945 86.680 ;
        RECT 102.230 86.520 102.400 87.490 ;
        RECT 102.685 87.330 102.855 89.860 ;
        RECT 103.275 89.840 103.445 89.860 ;
        RECT 103.730 89.655 103.900 91.065 ;
        RECT 104.185 90.860 104.355 90.880 ;
        RECT 104.775 90.860 104.945 90.880 ;
        RECT 104.155 90.445 104.385 90.860 ;
        RECT 104.745 90.445 104.975 90.860 ;
        RECT 104.155 90.275 104.975 90.445 ;
        RECT 104.155 89.860 104.385 90.275 ;
        RECT 104.745 89.860 104.975 90.275 ;
        RECT 104.185 89.840 104.355 89.860 ;
        RECT 104.775 89.840 104.945 89.860 ;
        RECT 105.230 89.655 105.400 91.065 ;
        RECT 105.685 90.860 105.855 90.880 ;
        RECT 106.275 90.860 106.445 91.455 ;
        RECT 106.585 91.065 107.045 91.295 ;
        RECT 105.655 89.860 105.885 90.860 ;
        RECT 106.245 89.860 106.475 90.860 ;
        RECT 103.585 89.425 104.045 89.655 ;
        RECT 105.085 89.425 105.545 89.655 ;
        RECT 103.730 87.720 103.900 89.425 ;
        RECT 104.110 88.465 104.430 88.725 ;
        RECT 103.585 87.490 104.045 87.720 ;
        RECT 103.275 87.330 103.445 87.350 ;
        RECT 102.655 86.680 102.885 87.330 ;
        RECT 103.245 86.680 103.475 87.330 ;
        RECT 102.685 86.660 102.855 86.680 ;
        RECT 102.085 86.290 102.545 86.520 ;
        RECT 103.275 86.085 103.445 86.680 ;
        RECT 103.730 86.565 103.900 87.490 ;
        RECT 104.185 87.330 104.355 88.465 ;
        RECT 105.230 87.720 105.400 89.425 ;
        RECT 105.685 88.725 105.855 89.860 ;
        RECT 106.275 89.840 106.445 89.860 ;
        RECT 106.730 89.655 106.900 91.065 ;
        RECT 107.140 90.635 107.400 90.955 ;
        RECT 107.155 89.860 107.385 90.635 ;
        RECT 106.585 89.425 107.045 89.655 ;
        RECT 106.730 88.725 106.900 89.425 ;
        RECT 105.610 88.465 105.930 88.725 ;
        RECT 106.655 88.465 106.975 88.725 ;
        RECT 105.085 87.490 105.545 87.720 ;
        RECT 104.775 87.330 104.945 87.350 ;
        RECT 104.155 86.680 104.385 87.330 ;
        RECT 104.745 86.680 104.975 87.330 ;
        RECT 104.185 86.660 104.355 86.680 ;
        RECT 103.685 86.520 103.945 86.565 ;
        RECT 103.585 86.290 104.045 86.520 ;
        RECT 103.685 86.245 103.945 86.290 ;
        RECT 104.775 86.085 104.945 86.680 ;
        RECT 105.230 86.565 105.400 87.490 ;
        RECT 105.685 87.330 105.855 88.465 ;
        RECT 106.730 87.720 106.900 88.465 ;
        RECT 106.585 87.490 107.045 87.720 ;
        RECT 106.275 87.330 106.445 87.350 ;
        RECT 105.655 86.680 105.885 87.330 ;
        RECT 106.245 86.680 106.475 87.330 ;
        RECT 105.685 86.660 105.855 86.680 ;
        RECT 105.185 86.520 105.445 86.565 ;
        RECT 105.085 86.290 105.545 86.520 ;
        RECT 105.185 86.245 105.445 86.290 ;
        RECT 105.185 86.085 105.445 86.100 ;
        RECT 106.275 86.085 106.445 86.680 ;
        RECT 106.730 86.520 106.900 87.490 ;
        RECT 107.185 87.330 107.355 89.860 ;
        RECT 107.670 89.440 107.990 91.280 ;
        RECT 107.155 86.680 107.385 87.330 ;
        RECT 107.185 86.660 107.355 86.680 ;
        RECT 106.585 86.290 107.045 86.520 ;
        RECT 31.065 85.795 107.565 86.085 ;
        RECT 31.685 85.780 31.945 85.795 ;
        RECT 105.185 85.780 105.445 85.795 ;
        RECT 33.185 85.400 33.445 85.475 ;
        RECT 36.185 85.400 36.445 85.475 ;
        RECT 83.325 85.400 83.585 85.475 ;
        RECT 33.185 85.230 83.585 85.400 ;
        RECT 33.185 85.155 33.445 85.230 ;
        RECT 36.185 85.155 36.445 85.230 ;
        RECT 83.325 85.155 83.585 85.230 ;
        RECT 37.685 85.015 37.945 85.090 ;
        RECT 40.685 85.015 40.945 85.090 ;
        RECT 86.310 85.015 86.570 85.090 ;
        RECT 37.685 84.845 86.570 85.015 ;
        RECT 37.685 84.770 37.945 84.845 ;
        RECT 40.685 84.770 40.945 84.845 ;
        RECT 86.310 84.770 86.570 84.845 ;
        RECT 34.820 84.695 35.120 84.725 ;
        RECT 30.550 84.395 35.120 84.695 ;
        RECT 34.820 84.365 35.120 84.395 ;
        RECT 42.185 84.630 42.445 84.705 ;
        RECT 45.185 84.630 45.445 84.705 ;
        RECT 76.115 84.630 76.375 84.705 ;
        RECT 42.185 84.460 76.375 84.630 ;
        RECT 42.185 84.385 42.445 84.460 ;
        RECT 45.185 84.385 45.445 84.460 ;
        RECT 76.115 84.385 76.375 84.460 ;
        RECT 105.360 84.695 105.660 84.725 ;
        RECT 107.830 84.695 108.130 87.740 ;
        RECT 105.360 84.395 108.130 84.695 ;
        RECT 105.360 84.365 105.660 84.395 ;
        RECT 46.685 84.245 46.945 84.320 ;
        RECT 49.685 84.245 49.945 84.320 ;
        RECT 79.600 84.245 79.860 84.320 ;
        RECT 46.685 84.075 79.860 84.245 ;
        RECT 46.685 84.000 46.945 84.075 ;
        RECT 49.685 84.000 49.945 84.075 ;
        RECT 79.600 84.000 79.860 84.075 ;
        RECT 51.185 83.860 51.445 83.935 ;
        RECT 54.185 83.860 54.445 83.935 ;
        RECT 69.905 83.860 70.165 83.935 ;
        RECT 51.185 83.690 70.165 83.860 ;
        RECT 51.185 83.615 51.445 83.690 ;
        RECT 54.185 83.615 54.445 83.690 ;
        RECT 69.905 83.615 70.165 83.690 ;
        RECT 55.685 83.475 55.945 83.550 ;
        RECT 58.685 83.475 58.945 83.550 ;
        RECT 72.890 83.475 73.150 83.550 ;
        RECT 55.685 83.305 73.150 83.475 ;
        RECT 55.685 83.230 55.945 83.305 ;
        RECT 58.685 83.230 58.945 83.305 ;
        RECT 72.890 83.230 73.150 83.305 ;
        RECT 60.185 83.090 60.445 83.165 ;
        RECT 62.695 83.090 62.955 83.165 ;
        RECT 63.185 83.090 63.445 83.165 ;
        RECT 60.185 82.920 63.445 83.090 ;
        RECT 60.185 82.845 60.445 82.920 ;
        RECT 62.695 82.845 62.955 82.920 ;
        RECT 63.185 82.845 63.445 82.920 ;
        RECT 64.685 82.705 64.945 82.780 ;
        RECT 66.180 82.705 66.440 82.780 ;
        RECT 67.685 82.705 67.945 82.780 ;
        RECT 64.685 82.535 67.945 82.705 ;
        RECT 64.685 82.460 64.945 82.535 ;
        RECT 66.180 82.460 66.440 82.535 ;
        RECT 67.685 82.460 67.945 82.535 ;
        RECT 55.985 82.320 56.245 82.395 ;
        RECT 69.185 82.320 69.445 82.395 ;
        RECT 72.185 82.320 72.445 82.395 ;
        RECT 55.985 82.150 72.445 82.320 ;
        RECT 55.985 82.075 56.245 82.150 ;
        RECT 69.185 82.075 69.445 82.150 ;
        RECT 72.185 82.075 72.445 82.150 ;
        RECT 59.470 81.935 59.730 82.010 ;
        RECT 73.685 81.935 73.945 82.010 ;
        RECT 76.685 81.935 76.945 82.010 ;
        RECT 59.470 81.765 76.945 81.935 ;
        RECT 59.470 81.690 59.730 81.765 ;
        RECT 73.685 81.690 73.945 81.765 ;
        RECT 76.685 81.690 76.945 81.765 ;
        RECT 49.275 81.550 49.535 81.625 ;
        RECT 78.185 81.550 78.445 81.625 ;
        RECT 81.185 81.550 81.445 81.625 ;
        RECT 49.275 81.380 81.445 81.550 ;
        RECT 49.275 81.305 49.535 81.380 ;
        RECT 78.185 81.305 78.445 81.380 ;
        RECT 81.185 81.305 81.445 81.380 ;
        RECT 52.760 81.165 53.020 81.240 ;
        RECT 82.685 81.165 82.945 81.240 ;
        RECT 85.685 81.165 85.945 81.240 ;
        RECT 52.760 80.995 85.945 81.165 ;
        RECT 52.760 80.920 53.020 80.995 ;
        RECT 82.685 80.920 82.945 80.995 ;
        RECT 85.685 80.920 85.945 80.995 ;
        RECT 42.565 80.780 42.825 80.855 ;
        RECT 87.185 80.780 87.445 80.855 ;
        RECT 90.185 80.780 90.445 80.855 ;
        RECT 42.565 80.610 90.445 80.780 ;
        RECT 42.565 80.535 42.825 80.610 ;
        RECT 87.185 80.535 87.445 80.610 ;
        RECT 90.185 80.535 90.445 80.610 ;
        RECT 46.050 80.395 46.310 80.470 ;
        RECT 91.685 80.395 91.945 80.470 ;
        RECT 94.685 80.395 94.945 80.470 ;
        RECT 46.050 80.225 94.945 80.395 ;
        RECT 46.050 80.150 46.310 80.225 ;
        RECT 91.685 80.150 91.945 80.225 ;
        RECT 94.685 80.150 94.945 80.225 ;
        RECT 35.855 80.010 36.115 80.085 ;
        RECT 96.185 80.010 96.445 80.085 ;
        RECT 99.185 80.010 99.445 80.085 ;
        RECT 35.855 79.840 99.445 80.010 ;
        RECT 35.855 79.765 36.115 79.840 ;
        RECT 96.185 79.765 96.445 79.840 ;
        RECT 99.185 79.765 99.445 79.840 ;
        RECT 39.340 79.625 39.600 79.700 ;
        RECT 100.685 79.625 100.945 79.700 ;
        RECT 103.685 79.625 103.945 79.700 ;
        RECT 39.340 79.455 103.945 79.625 ;
        RECT 39.340 79.380 39.600 79.455 ;
        RECT 100.685 79.380 100.945 79.455 ;
        RECT 103.685 79.380 103.945 79.455 ;
        RECT 36.320 77.635 36.610 78.500 ;
        RECT 37.205 78.290 38.205 78.320 ;
        RECT 39.340 78.290 39.600 78.365 ;
        RECT 40.735 78.290 41.385 78.320 ;
        RECT 37.185 78.120 41.405 78.290 ;
        RECT 37.205 78.090 38.205 78.120 ;
        RECT 39.340 78.045 39.600 78.120 ;
        RECT 40.735 78.090 41.385 78.120 ;
        RECT 36.770 77.835 37.000 77.980 ;
        RECT 37.185 77.835 37.445 77.910 ;
        RECT 38.410 77.835 38.640 77.980 ;
        RECT 40.345 77.835 40.575 77.980 ;
        RECT 41.545 77.835 41.775 77.980 ;
        RECT 36.770 77.665 41.775 77.835 ;
        RECT 36.315 77.275 36.615 77.635 ;
        RECT 36.770 77.520 37.000 77.665 ;
        RECT 37.185 77.590 37.445 77.665 ;
        RECT 38.410 77.520 38.640 77.665 ;
        RECT 40.345 77.520 40.575 77.665 ;
        RECT 41.545 77.520 41.775 77.665 ;
        RECT 37.205 77.380 38.205 77.410 ;
        RECT 40.735 77.380 41.385 77.410 ;
        RECT 41.980 77.380 42.270 78.500 ;
        RECT 43.030 77.635 43.320 78.500 ;
        RECT 43.915 78.290 44.915 78.320 ;
        RECT 46.050 78.290 46.310 78.365 ;
        RECT 47.445 78.290 48.095 78.320 ;
        RECT 43.895 78.120 48.115 78.290 ;
        RECT 43.915 78.090 44.915 78.120 ;
        RECT 46.050 78.045 46.310 78.120 ;
        RECT 47.445 78.090 48.095 78.120 ;
        RECT 43.480 77.835 43.710 77.980 ;
        RECT 43.895 77.835 44.155 77.910 ;
        RECT 45.120 77.835 45.350 77.980 ;
        RECT 47.055 77.835 47.285 77.980 ;
        RECT 48.255 77.835 48.485 77.980 ;
        RECT 43.480 77.665 48.485 77.835 ;
        RECT 36.320 74.635 36.610 77.275 ;
        RECT 37.185 77.210 38.225 77.380 ;
        RECT 40.715 77.210 42.270 77.380 ;
        RECT 43.025 77.275 43.325 77.635 ;
        RECT 43.480 77.520 43.710 77.665 ;
        RECT 43.895 77.590 44.155 77.665 ;
        RECT 45.120 77.520 45.350 77.665 ;
        RECT 47.055 77.520 47.285 77.665 ;
        RECT 48.255 77.520 48.485 77.665 ;
        RECT 43.915 77.380 44.915 77.410 ;
        RECT 47.445 77.380 48.095 77.410 ;
        RECT 48.690 77.380 48.980 78.500 ;
        RECT 49.740 77.635 50.030 78.500 ;
        RECT 50.625 78.290 51.625 78.320 ;
        RECT 52.760 78.290 53.020 78.365 ;
        RECT 54.155 78.290 54.805 78.320 ;
        RECT 50.605 78.120 54.825 78.290 ;
        RECT 50.625 78.090 51.625 78.120 ;
        RECT 52.760 78.045 53.020 78.120 ;
        RECT 54.155 78.090 54.805 78.120 ;
        RECT 50.190 77.835 50.420 77.980 ;
        RECT 50.605 77.835 50.865 77.910 ;
        RECT 51.830 77.835 52.060 77.980 ;
        RECT 53.765 77.835 53.995 77.980 ;
        RECT 54.965 77.835 55.195 77.980 ;
        RECT 50.190 77.665 55.195 77.835 ;
        RECT 37.205 77.180 38.205 77.210 ;
        RECT 40.735 77.180 41.385 77.210 ;
        RECT 37.620 76.820 37.790 77.180 ;
        RECT 37.205 76.790 38.205 76.820 ;
        RECT 39.340 76.790 39.600 76.865 ;
        RECT 40.735 76.790 41.385 76.820 ;
        RECT 37.185 76.620 38.225 76.790 ;
        RECT 39.340 76.620 41.405 76.790 ;
        RECT 37.205 76.590 38.205 76.620 ;
        RECT 39.340 76.545 39.600 76.620 ;
        RECT 40.735 76.590 41.385 76.620 ;
        RECT 36.770 76.335 37.000 76.480 ;
        RECT 38.410 76.410 38.640 76.480 ;
        RECT 38.025 76.335 38.640 76.410 ;
        RECT 40.345 76.335 40.575 76.480 ;
        RECT 41.545 76.335 41.775 76.480 ;
        RECT 36.770 76.165 41.775 76.335 ;
        RECT 36.770 76.020 37.000 76.165 ;
        RECT 38.025 76.090 38.640 76.165 ;
        RECT 38.410 76.020 38.640 76.090 ;
        RECT 40.345 76.020 40.575 76.165 ;
        RECT 41.545 76.020 41.775 76.165 ;
        RECT 41.980 76.135 42.270 77.210 ;
        RECT 37.205 75.880 38.205 75.910 ;
        RECT 40.735 75.880 41.385 75.910 ;
        RECT 41.975 75.880 42.275 76.135 ;
        RECT 37.185 75.710 38.225 75.880 ;
        RECT 40.715 75.775 42.275 75.880 ;
        RECT 40.715 75.710 42.270 75.775 ;
        RECT 37.205 75.680 38.205 75.710 ;
        RECT 40.735 75.680 41.385 75.710 ;
        RECT 37.620 75.320 37.790 75.680 ;
        RECT 37.205 75.290 38.205 75.320 ;
        RECT 39.340 75.290 39.600 75.365 ;
        RECT 40.735 75.290 41.385 75.320 ;
        RECT 37.185 75.120 38.225 75.290 ;
        RECT 39.340 75.120 41.405 75.290 ;
        RECT 37.205 75.090 38.205 75.120 ;
        RECT 39.340 75.045 39.600 75.120 ;
        RECT 40.735 75.090 41.385 75.120 ;
        RECT 36.770 74.835 37.000 74.980 ;
        RECT 38.410 74.910 38.640 74.980 ;
        RECT 38.410 74.835 38.705 74.910 ;
        RECT 40.345 74.835 40.575 74.980 ;
        RECT 41.545 74.835 41.775 74.980 ;
        RECT 36.770 74.665 41.775 74.835 ;
        RECT 36.315 74.380 36.615 74.635 ;
        RECT 36.770 74.520 37.000 74.665 ;
        RECT 38.410 74.590 38.705 74.665 ;
        RECT 38.410 74.520 38.640 74.590 ;
        RECT 40.345 74.520 40.575 74.665 ;
        RECT 41.545 74.520 41.775 74.665 ;
        RECT 37.205 74.380 38.205 74.410 ;
        RECT 40.735 74.380 41.385 74.410 ;
        RECT 41.980 74.380 42.270 75.710 ;
        RECT 43.030 74.635 43.320 77.275 ;
        RECT 43.895 77.210 44.935 77.380 ;
        RECT 47.425 77.210 48.980 77.380 ;
        RECT 49.735 77.275 50.035 77.635 ;
        RECT 50.190 77.520 50.420 77.665 ;
        RECT 50.605 77.590 50.865 77.665 ;
        RECT 51.830 77.520 52.060 77.665 ;
        RECT 53.765 77.520 53.995 77.665 ;
        RECT 54.965 77.520 55.195 77.665 ;
        RECT 50.625 77.380 51.625 77.410 ;
        RECT 54.155 77.380 54.805 77.410 ;
        RECT 55.400 77.380 55.690 78.500 ;
        RECT 56.450 77.635 56.740 78.500 ;
        RECT 57.335 78.290 58.335 78.320 ;
        RECT 59.470 78.290 59.730 78.365 ;
        RECT 60.865 78.290 61.515 78.320 ;
        RECT 57.315 78.120 61.535 78.290 ;
        RECT 57.335 78.090 58.335 78.120 ;
        RECT 59.470 78.045 59.730 78.120 ;
        RECT 60.865 78.090 61.515 78.120 ;
        RECT 56.900 77.835 57.130 77.980 ;
        RECT 57.315 77.835 57.575 77.910 ;
        RECT 58.540 77.835 58.770 77.980 ;
        RECT 60.475 77.835 60.705 77.980 ;
        RECT 61.675 77.835 61.905 77.980 ;
        RECT 56.900 77.665 61.905 77.835 ;
        RECT 43.915 77.180 44.915 77.210 ;
        RECT 47.445 77.180 48.095 77.210 ;
        RECT 44.330 76.820 44.500 77.180 ;
        RECT 43.915 76.790 44.915 76.820 ;
        RECT 46.050 76.790 46.310 76.865 ;
        RECT 47.445 76.790 48.095 76.820 ;
        RECT 43.895 76.620 44.935 76.790 ;
        RECT 46.050 76.620 48.115 76.790 ;
        RECT 43.915 76.590 44.915 76.620 ;
        RECT 46.050 76.545 46.310 76.620 ;
        RECT 47.445 76.590 48.095 76.620 ;
        RECT 43.480 76.335 43.710 76.480 ;
        RECT 45.120 76.410 45.350 76.480 ;
        RECT 44.735 76.335 45.350 76.410 ;
        RECT 47.055 76.335 47.285 76.480 ;
        RECT 48.255 76.335 48.485 76.480 ;
        RECT 43.480 76.165 48.485 76.335 ;
        RECT 43.480 76.020 43.710 76.165 ;
        RECT 44.735 76.090 45.350 76.165 ;
        RECT 45.120 76.020 45.350 76.090 ;
        RECT 47.055 76.020 47.285 76.165 ;
        RECT 48.255 76.020 48.485 76.165 ;
        RECT 48.690 76.135 48.980 77.210 ;
        RECT 43.915 75.880 44.915 75.910 ;
        RECT 47.445 75.880 48.095 75.910 ;
        RECT 48.685 75.880 48.985 76.135 ;
        RECT 43.895 75.710 44.935 75.880 ;
        RECT 47.425 75.775 48.985 75.880 ;
        RECT 47.425 75.710 48.980 75.775 ;
        RECT 43.915 75.680 44.915 75.710 ;
        RECT 47.445 75.680 48.095 75.710 ;
        RECT 44.330 75.320 44.500 75.680 ;
        RECT 43.915 75.290 44.915 75.320 ;
        RECT 46.050 75.290 46.310 75.365 ;
        RECT 47.445 75.290 48.095 75.320 ;
        RECT 43.895 75.120 44.935 75.290 ;
        RECT 46.050 75.120 48.115 75.290 ;
        RECT 43.915 75.090 44.915 75.120 ;
        RECT 46.050 75.045 46.310 75.120 ;
        RECT 47.445 75.090 48.095 75.120 ;
        RECT 43.480 74.835 43.710 74.980 ;
        RECT 45.120 74.910 45.350 74.980 ;
        RECT 45.120 74.835 45.415 74.910 ;
        RECT 47.055 74.835 47.285 74.980 ;
        RECT 48.255 74.835 48.485 74.980 ;
        RECT 43.480 74.665 48.485 74.835 ;
        RECT 36.315 74.275 38.225 74.380 ;
        RECT 36.320 74.210 38.225 74.275 ;
        RECT 40.715 74.210 42.270 74.380 ;
        RECT 43.025 74.380 43.325 74.635 ;
        RECT 43.480 74.520 43.710 74.665 ;
        RECT 45.120 74.590 45.415 74.665 ;
        RECT 45.120 74.520 45.350 74.590 ;
        RECT 47.055 74.520 47.285 74.665 ;
        RECT 48.255 74.520 48.485 74.665 ;
        RECT 43.915 74.380 44.915 74.410 ;
        RECT 47.445 74.380 48.095 74.410 ;
        RECT 48.690 74.380 48.980 75.710 ;
        RECT 49.740 74.635 50.030 77.275 ;
        RECT 50.605 77.210 51.645 77.380 ;
        RECT 54.135 77.210 55.690 77.380 ;
        RECT 56.445 77.275 56.745 77.635 ;
        RECT 56.900 77.520 57.130 77.665 ;
        RECT 57.315 77.590 57.575 77.665 ;
        RECT 58.540 77.520 58.770 77.665 ;
        RECT 60.475 77.520 60.705 77.665 ;
        RECT 61.675 77.520 61.905 77.665 ;
        RECT 57.335 77.380 58.335 77.410 ;
        RECT 60.865 77.380 61.515 77.410 ;
        RECT 62.110 77.380 62.400 78.500 ;
        RECT 63.160 77.635 63.450 78.500 ;
        RECT 64.045 78.290 65.045 78.320 ;
        RECT 66.180 78.290 66.440 78.365 ;
        RECT 67.575 78.290 68.225 78.320 ;
        RECT 64.025 78.120 68.245 78.290 ;
        RECT 64.045 78.090 65.045 78.120 ;
        RECT 66.180 78.045 66.440 78.120 ;
        RECT 67.575 78.090 68.225 78.120 ;
        RECT 63.610 77.835 63.840 77.980 ;
        RECT 64.025 77.835 64.285 77.910 ;
        RECT 65.250 77.835 65.480 77.980 ;
        RECT 67.185 77.835 67.415 77.980 ;
        RECT 68.385 77.835 68.615 77.980 ;
        RECT 63.610 77.665 68.615 77.835 ;
        RECT 50.625 77.180 51.625 77.210 ;
        RECT 54.155 77.180 54.805 77.210 ;
        RECT 51.040 76.820 51.210 77.180 ;
        RECT 50.625 76.790 51.625 76.820 ;
        RECT 52.760 76.790 53.020 76.865 ;
        RECT 54.155 76.790 54.805 76.820 ;
        RECT 50.605 76.620 51.645 76.790 ;
        RECT 52.760 76.620 54.825 76.790 ;
        RECT 50.625 76.590 51.625 76.620 ;
        RECT 52.760 76.545 53.020 76.620 ;
        RECT 54.155 76.590 54.805 76.620 ;
        RECT 50.190 76.335 50.420 76.480 ;
        RECT 51.830 76.410 52.060 76.480 ;
        RECT 51.445 76.335 52.060 76.410 ;
        RECT 53.765 76.335 53.995 76.480 ;
        RECT 54.965 76.335 55.195 76.480 ;
        RECT 50.190 76.165 55.195 76.335 ;
        RECT 50.190 76.020 50.420 76.165 ;
        RECT 51.445 76.090 52.060 76.165 ;
        RECT 51.830 76.020 52.060 76.090 ;
        RECT 53.765 76.020 53.995 76.165 ;
        RECT 54.965 76.020 55.195 76.165 ;
        RECT 55.400 76.135 55.690 77.210 ;
        RECT 50.625 75.880 51.625 75.910 ;
        RECT 54.155 75.880 54.805 75.910 ;
        RECT 55.395 75.880 55.695 76.135 ;
        RECT 50.605 75.710 51.645 75.880 ;
        RECT 54.135 75.775 55.695 75.880 ;
        RECT 54.135 75.710 55.690 75.775 ;
        RECT 50.625 75.680 51.625 75.710 ;
        RECT 54.155 75.680 54.805 75.710 ;
        RECT 51.040 75.320 51.210 75.680 ;
        RECT 50.625 75.290 51.625 75.320 ;
        RECT 52.760 75.290 53.020 75.365 ;
        RECT 54.155 75.290 54.805 75.320 ;
        RECT 50.605 75.120 51.645 75.290 ;
        RECT 52.760 75.120 54.825 75.290 ;
        RECT 50.625 75.090 51.625 75.120 ;
        RECT 52.760 75.045 53.020 75.120 ;
        RECT 54.155 75.090 54.805 75.120 ;
        RECT 50.190 74.835 50.420 74.980 ;
        RECT 51.830 74.910 52.060 74.980 ;
        RECT 51.830 74.835 52.125 74.910 ;
        RECT 53.765 74.835 53.995 74.980 ;
        RECT 54.965 74.835 55.195 74.980 ;
        RECT 50.190 74.665 55.195 74.835 ;
        RECT 43.025 74.275 44.935 74.380 ;
        RECT 36.320 71.635 36.610 74.210 ;
        RECT 37.205 74.180 38.205 74.210 ;
        RECT 40.735 74.180 41.385 74.210 ;
        RECT 37.205 73.790 38.205 73.820 ;
        RECT 39.340 73.790 39.600 73.865 ;
        RECT 40.735 73.790 41.385 73.820 ;
        RECT 37.185 73.620 41.405 73.790 ;
        RECT 37.205 73.590 38.205 73.620 ;
        RECT 39.340 73.545 39.600 73.620 ;
        RECT 40.735 73.590 41.385 73.620 ;
        RECT 36.770 73.335 37.000 73.480 ;
        RECT 37.185 73.335 37.445 73.410 ;
        RECT 38.410 73.335 38.640 73.480 ;
        RECT 40.345 73.335 40.575 73.480 ;
        RECT 41.545 73.335 41.775 73.480 ;
        RECT 36.770 73.165 41.775 73.335 ;
        RECT 36.770 73.020 37.000 73.165 ;
        RECT 37.185 73.090 37.445 73.165 ;
        RECT 38.410 73.020 38.640 73.165 ;
        RECT 40.345 73.020 40.575 73.165 ;
        RECT 41.545 73.020 41.775 73.165 ;
        RECT 41.980 73.135 42.270 74.210 ;
        RECT 43.030 74.210 44.935 74.275 ;
        RECT 47.425 74.210 48.980 74.380 ;
        RECT 49.735 74.380 50.035 74.635 ;
        RECT 50.190 74.520 50.420 74.665 ;
        RECT 51.830 74.590 52.125 74.665 ;
        RECT 51.830 74.520 52.060 74.590 ;
        RECT 53.765 74.520 53.995 74.665 ;
        RECT 54.965 74.520 55.195 74.665 ;
        RECT 50.625 74.380 51.625 74.410 ;
        RECT 54.155 74.380 54.805 74.410 ;
        RECT 55.400 74.380 55.690 75.710 ;
        RECT 56.450 74.635 56.740 77.275 ;
        RECT 57.315 77.210 58.355 77.380 ;
        RECT 60.845 77.210 62.400 77.380 ;
        RECT 63.155 77.275 63.455 77.635 ;
        RECT 63.610 77.520 63.840 77.665 ;
        RECT 64.025 77.590 64.285 77.665 ;
        RECT 65.250 77.520 65.480 77.665 ;
        RECT 67.185 77.520 67.415 77.665 ;
        RECT 68.385 77.520 68.615 77.665 ;
        RECT 64.045 77.380 65.045 77.410 ;
        RECT 67.575 77.380 68.225 77.410 ;
        RECT 68.820 77.380 69.110 78.500 ;
        RECT 69.870 77.635 70.160 78.500 ;
        RECT 70.755 78.290 71.755 78.320 ;
        RECT 72.890 78.290 73.150 78.365 ;
        RECT 74.285 78.290 74.935 78.320 ;
        RECT 70.735 78.120 74.955 78.290 ;
        RECT 70.755 78.090 71.755 78.120 ;
        RECT 72.890 78.045 73.150 78.120 ;
        RECT 74.285 78.090 74.935 78.120 ;
        RECT 70.320 77.835 70.550 77.980 ;
        RECT 70.735 77.835 70.995 77.910 ;
        RECT 71.960 77.835 72.190 77.980 ;
        RECT 73.895 77.835 74.125 77.980 ;
        RECT 75.095 77.835 75.325 77.980 ;
        RECT 70.320 77.665 75.325 77.835 ;
        RECT 57.335 77.180 58.335 77.210 ;
        RECT 60.865 77.180 61.515 77.210 ;
        RECT 57.750 76.820 57.920 77.180 ;
        RECT 57.335 76.790 58.335 76.820 ;
        RECT 59.470 76.790 59.730 76.865 ;
        RECT 60.865 76.790 61.515 76.820 ;
        RECT 57.315 76.620 58.355 76.790 ;
        RECT 59.470 76.620 61.535 76.790 ;
        RECT 57.335 76.590 58.335 76.620 ;
        RECT 59.470 76.545 59.730 76.620 ;
        RECT 60.865 76.590 61.515 76.620 ;
        RECT 56.900 76.335 57.130 76.480 ;
        RECT 58.540 76.410 58.770 76.480 ;
        RECT 58.155 76.335 58.770 76.410 ;
        RECT 60.475 76.335 60.705 76.480 ;
        RECT 61.675 76.335 61.905 76.480 ;
        RECT 56.900 76.165 61.905 76.335 ;
        RECT 56.900 76.020 57.130 76.165 ;
        RECT 58.155 76.090 58.770 76.165 ;
        RECT 58.540 76.020 58.770 76.090 ;
        RECT 60.475 76.020 60.705 76.165 ;
        RECT 61.675 76.020 61.905 76.165 ;
        RECT 62.110 76.135 62.400 77.210 ;
        RECT 57.335 75.880 58.335 75.910 ;
        RECT 60.865 75.880 61.515 75.910 ;
        RECT 62.105 75.880 62.405 76.135 ;
        RECT 57.315 75.710 58.355 75.880 ;
        RECT 60.845 75.775 62.405 75.880 ;
        RECT 60.845 75.710 62.400 75.775 ;
        RECT 57.335 75.680 58.335 75.710 ;
        RECT 60.865 75.680 61.515 75.710 ;
        RECT 57.750 75.320 57.920 75.680 ;
        RECT 57.335 75.290 58.335 75.320 ;
        RECT 59.470 75.290 59.730 75.365 ;
        RECT 60.865 75.290 61.515 75.320 ;
        RECT 57.315 75.120 58.355 75.290 ;
        RECT 59.470 75.120 61.535 75.290 ;
        RECT 57.335 75.090 58.335 75.120 ;
        RECT 59.470 75.045 59.730 75.120 ;
        RECT 60.865 75.090 61.515 75.120 ;
        RECT 56.900 74.835 57.130 74.980 ;
        RECT 58.540 74.910 58.770 74.980 ;
        RECT 58.540 74.835 58.835 74.910 ;
        RECT 60.475 74.835 60.705 74.980 ;
        RECT 61.675 74.835 61.905 74.980 ;
        RECT 56.900 74.665 61.905 74.835 ;
        RECT 49.735 74.275 51.645 74.380 ;
        RECT 37.205 72.880 38.205 72.910 ;
        RECT 40.735 72.880 41.385 72.910 ;
        RECT 41.975 72.880 42.275 73.135 ;
        RECT 37.185 72.710 38.225 72.880 ;
        RECT 40.715 72.775 42.275 72.880 ;
        RECT 40.715 72.710 42.270 72.775 ;
        RECT 37.205 72.680 38.205 72.710 ;
        RECT 40.735 72.680 41.385 72.710 ;
        RECT 37.620 72.320 37.790 72.680 ;
        RECT 37.205 72.290 38.205 72.320 ;
        RECT 39.340 72.290 39.600 72.365 ;
        RECT 40.735 72.290 41.385 72.320 ;
        RECT 37.185 72.120 38.225 72.290 ;
        RECT 39.340 72.120 41.405 72.290 ;
        RECT 37.205 72.090 38.205 72.120 ;
        RECT 39.340 72.045 39.600 72.120 ;
        RECT 40.735 72.090 41.385 72.120 ;
        RECT 36.770 71.835 37.000 71.980 ;
        RECT 37.605 71.835 37.865 71.910 ;
        RECT 38.410 71.835 38.640 71.980 ;
        RECT 40.345 71.835 40.575 71.980 ;
        RECT 41.545 71.835 41.775 71.980 ;
        RECT 36.770 71.665 41.775 71.835 ;
        RECT 36.315 71.275 36.615 71.635 ;
        RECT 36.770 71.520 37.000 71.665 ;
        RECT 37.605 71.590 37.865 71.665 ;
        RECT 38.410 71.520 38.640 71.665 ;
        RECT 40.345 71.520 40.575 71.665 ;
        RECT 41.545 71.520 41.775 71.665 ;
        RECT 37.205 71.380 38.205 71.410 ;
        RECT 40.735 71.380 41.385 71.410 ;
        RECT 41.980 71.380 42.270 72.710 ;
        RECT 43.030 71.635 43.320 74.210 ;
        RECT 43.915 74.180 44.915 74.210 ;
        RECT 47.445 74.180 48.095 74.210 ;
        RECT 43.915 73.790 44.915 73.820 ;
        RECT 46.050 73.790 46.310 73.865 ;
        RECT 47.445 73.790 48.095 73.820 ;
        RECT 43.895 73.620 48.115 73.790 ;
        RECT 43.915 73.590 44.915 73.620 ;
        RECT 46.050 73.545 46.310 73.620 ;
        RECT 47.445 73.590 48.095 73.620 ;
        RECT 43.480 73.335 43.710 73.480 ;
        RECT 43.895 73.335 44.155 73.410 ;
        RECT 45.120 73.335 45.350 73.480 ;
        RECT 47.055 73.335 47.285 73.480 ;
        RECT 48.255 73.335 48.485 73.480 ;
        RECT 43.480 73.165 48.485 73.335 ;
        RECT 43.480 73.020 43.710 73.165 ;
        RECT 43.895 73.090 44.155 73.165 ;
        RECT 45.120 73.020 45.350 73.165 ;
        RECT 47.055 73.020 47.285 73.165 ;
        RECT 48.255 73.020 48.485 73.165 ;
        RECT 48.690 73.135 48.980 74.210 ;
        RECT 49.740 74.210 51.645 74.275 ;
        RECT 54.135 74.210 55.690 74.380 ;
        RECT 56.445 74.380 56.745 74.635 ;
        RECT 56.900 74.520 57.130 74.665 ;
        RECT 58.540 74.590 58.835 74.665 ;
        RECT 58.540 74.520 58.770 74.590 ;
        RECT 60.475 74.520 60.705 74.665 ;
        RECT 61.675 74.520 61.905 74.665 ;
        RECT 57.335 74.380 58.335 74.410 ;
        RECT 60.865 74.380 61.515 74.410 ;
        RECT 62.110 74.380 62.400 75.710 ;
        RECT 63.160 74.635 63.450 77.275 ;
        RECT 64.025 77.210 65.065 77.380 ;
        RECT 67.555 77.210 69.110 77.380 ;
        RECT 69.865 77.275 70.165 77.635 ;
        RECT 70.320 77.520 70.550 77.665 ;
        RECT 70.735 77.590 70.995 77.665 ;
        RECT 71.960 77.520 72.190 77.665 ;
        RECT 73.895 77.520 74.125 77.665 ;
        RECT 75.095 77.520 75.325 77.665 ;
        RECT 70.755 77.380 71.755 77.410 ;
        RECT 74.285 77.380 74.935 77.410 ;
        RECT 75.530 77.380 75.820 78.500 ;
        RECT 76.580 77.635 76.870 78.500 ;
        RECT 77.465 78.290 78.465 78.320 ;
        RECT 79.600 78.290 79.860 78.365 ;
        RECT 80.995 78.290 81.645 78.320 ;
        RECT 77.445 78.120 81.665 78.290 ;
        RECT 77.465 78.090 78.465 78.120 ;
        RECT 79.600 78.045 79.860 78.120 ;
        RECT 80.995 78.090 81.645 78.120 ;
        RECT 77.030 77.835 77.260 77.980 ;
        RECT 77.445 77.835 77.705 77.910 ;
        RECT 78.670 77.835 78.900 77.980 ;
        RECT 80.605 77.835 80.835 77.980 ;
        RECT 81.805 77.835 82.035 77.980 ;
        RECT 77.030 77.665 82.035 77.835 ;
        RECT 64.045 77.180 65.045 77.210 ;
        RECT 67.575 77.180 68.225 77.210 ;
        RECT 64.460 76.820 64.630 77.180 ;
        RECT 64.045 76.790 65.045 76.820 ;
        RECT 66.180 76.790 66.440 76.865 ;
        RECT 67.575 76.790 68.225 76.820 ;
        RECT 64.025 76.620 65.065 76.790 ;
        RECT 66.180 76.620 68.245 76.790 ;
        RECT 64.045 76.590 65.045 76.620 ;
        RECT 66.180 76.545 66.440 76.620 ;
        RECT 67.575 76.590 68.225 76.620 ;
        RECT 63.610 76.335 63.840 76.480 ;
        RECT 65.250 76.410 65.480 76.480 ;
        RECT 64.865 76.335 65.480 76.410 ;
        RECT 67.185 76.335 67.415 76.480 ;
        RECT 68.385 76.335 68.615 76.480 ;
        RECT 63.610 76.165 68.615 76.335 ;
        RECT 63.610 76.020 63.840 76.165 ;
        RECT 64.865 76.090 65.480 76.165 ;
        RECT 65.250 76.020 65.480 76.090 ;
        RECT 67.185 76.020 67.415 76.165 ;
        RECT 68.385 76.020 68.615 76.165 ;
        RECT 68.820 76.135 69.110 77.210 ;
        RECT 64.045 75.880 65.045 75.910 ;
        RECT 67.575 75.880 68.225 75.910 ;
        RECT 68.815 75.880 69.115 76.135 ;
        RECT 64.025 75.710 65.065 75.880 ;
        RECT 67.555 75.775 69.115 75.880 ;
        RECT 67.555 75.710 69.110 75.775 ;
        RECT 64.045 75.680 65.045 75.710 ;
        RECT 67.575 75.680 68.225 75.710 ;
        RECT 64.460 75.320 64.630 75.680 ;
        RECT 64.045 75.290 65.045 75.320 ;
        RECT 66.180 75.290 66.440 75.365 ;
        RECT 67.575 75.290 68.225 75.320 ;
        RECT 64.025 75.120 65.065 75.290 ;
        RECT 66.180 75.120 68.245 75.290 ;
        RECT 64.045 75.090 65.045 75.120 ;
        RECT 66.180 75.045 66.440 75.120 ;
        RECT 67.575 75.090 68.225 75.120 ;
        RECT 63.610 74.835 63.840 74.980 ;
        RECT 65.250 74.910 65.480 74.980 ;
        RECT 65.250 74.835 65.545 74.910 ;
        RECT 67.185 74.835 67.415 74.980 ;
        RECT 68.385 74.835 68.615 74.980 ;
        RECT 63.610 74.665 68.615 74.835 ;
        RECT 56.445 74.275 58.355 74.380 ;
        RECT 43.915 72.880 44.915 72.910 ;
        RECT 47.445 72.880 48.095 72.910 ;
        RECT 48.685 72.880 48.985 73.135 ;
        RECT 43.895 72.710 44.935 72.880 ;
        RECT 47.425 72.775 48.985 72.880 ;
        RECT 47.425 72.710 48.980 72.775 ;
        RECT 43.915 72.680 44.915 72.710 ;
        RECT 47.445 72.680 48.095 72.710 ;
        RECT 44.330 72.320 44.500 72.680 ;
        RECT 43.915 72.290 44.915 72.320 ;
        RECT 46.050 72.290 46.310 72.365 ;
        RECT 47.445 72.290 48.095 72.320 ;
        RECT 43.895 72.120 44.935 72.290 ;
        RECT 46.050 72.120 48.115 72.290 ;
        RECT 43.915 72.090 44.915 72.120 ;
        RECT 46.050 72.045 46.310 72.120 ;
        RECT 47.445 72.090 48.095 72.120 ;
        RECT 43.480 71.835 43.710 71.980 ;
        RECT 44.315 71.835 44.575 71.910 ;
        RECT 45.120 71.835 45.350 71.980 ;
        RECT 47.055 71.835 47.285 71.980 ;
        RECT 48.255 71.835 48.485 71.980 ;
        RECT 43.480 71.665 48.485 71.835 ;
        RECT 36.320 69.880 36.610 71.275 ;
        RECT 37.185 71.210 38.225 71.380 ;
        RECT 40.715 71.210 42.270 71.380 ;
        RECT 43.025 71.275 43.325 71.635 ;
        RECT 43.480 71.520 43.710 71.665 ;
        RECT 44.315 71.590 44.575 71.665 ;
        RECT 45.120 71.520 45.350 71.665 ;
        RECT 47.055 71.520 47.285 71.665 ;
        RECT 48.255 71.520 48.485 71.665 ;
        RECT 43.915 71.380 44.915 71.410 ;
        RECT 47.445 71.380 48.095 71.410 ;
        RECT 48.690 71.380 48.980 72.710 ;
        RECT 49.740 71.635 50.030 74.210 ;
        RECT 50.625 74.180 51.625 74.210 ;
        RECT 54.155 74.180 54.805 74.210 ;
        RECT 50.625 73.790 51.625 73.820 ;
        RECT 52.760 73.790 53.020 73.865 ;
        RECT 54.155 73.790 54.805 73.820 ;
        RECT 50.605 73.620 54.825 73.790 ;
        RECT 50.625 73.590 51.625 73.620 ;
        RECT 52.760 73.545 53.020 73.620 ;
        RECT 54.155 73.590 54.805 73.620 ;
        RECT 50.190 73.335 50.420 73.480 ;
        RECT 50.605 73.335 50.865 73.410 ;
        RECT 51.830 73.335 52.060 73.480 ;
        RECT 53.765 73.335 53.995 73.480 ;
        RECT 54.965 73.335 55.195 73.480 ;
        RECT 50.190 73.165 55.195 73.335 ;
        RECT 50.190 73.020 50.420 73.165 ;
        RECT 50.605 73.090 50.865 73.165 ;
        RECT 51.830 73.020 52.060 73.165 ;
        RECT 53.765 73.020 53.995 73.165 ;
        RECT 54.965 73.020 55.195 73.165 ;
        RECT 55.400 73.135 55.690 74.210 ;
        RECT 56.450 74.210 58.355 74.275 ;
        RECT 60.845 74.210 62.400 74.380 ;
        RECT 63.155 74.380 63.455 74.635 ;
        RECT 63.610 74.520 63.840 74.665 ;
        RECT 65.250 74.590 65.545 74.665 ;
        RECT 65.250 74.520 65.480 74.590 ;
        RECT 67.185 74.520 67.415 74.665 ;
        RECT 68.385 74.520 68.615 74.665 ;
        RECT 64.045 74.380 65.045 74.410 ;
        RECT 67.575 74.380 68.225 74.410 ;
        RECT 68.820 74.380 69.110 75.710 ;
        RECT 69.870 74.635 70.160 77.275 ;
        RECT 70.735 77.210 71.775 77.380 ;
        RECT 74.265 77.210 75.820 77.380 ;
        RECT 76.575 77.275 76.875 77.635 ;
        RECT 77.030 77.520 77.260 77.665 ;
        RECT 77.445 77.590 77.705 77.665 ;
        RECT 78.670 77.520 78.900 77.665 ;
        RECT 80.605 77.520 80.835 77.665 ;
        RECT 81.805 77.520 82.035 77.665 ;
        RECT 77.465 77.380 78.465 77.410 ;
        RECT 80.995 77.380 81.645 77.410 ;
        RECT 82.240 77.380 82.530 78.500 ;
        RECT 83.290 77.635 83.580 78.500 ;
        RECT 84.175 78.290 85.175 78.320 ;
        RECT 86.310 78.290 86.570 78.365 ;
        RECT 87.705 78.290 88.355 78.320 ;
        RECT 84.155 78.120 88.375 78.290 ;
        RECT 84.175 78.090 85.175 78.120 ;
        RECT 86.310 78.045 86.570 78.120 ;
        RECT 87.705 78.090 88.355 78.120 ;
        RECT 83.740 77.835 83.970 77.980 ;
        RECT 84.155 77.835 84.415 77.910 ;
        RECT 85.380 77.835 85.610 77.980 ;
        RECT 87.315 77.835 87.545 77.980 ;
        RECT 88.515 77.835 88.745 77.980 ;
        RECT 83.740 77.665 88.745 77.835 ;
        RECT 70.755 77.180 71.755 77.210 ;
        RECT 74.285 77.180 74.935 77.210 ;
        RECT 71.170 76.820 71.340 77.180 ;
        RECT 70.755 76.790 71.755 76.820 ;
        RECT 72.890 76.790 73.150 76.865 ;
        RECT 74.285 76.790 74.935 76.820 ;
        RECT 70.735 76.620 71.775 76.790 ;
        RECT 72.890 76.620 74.955 76.790 ;
        RECT 70.755 76.590 71.755 76.620 ;
        RECT 72.890 76.545 73.150 76.620 ;
        RECT 74.285 76.590 74.935 76.620 ;
        RECT 70.320 76.335 70.550 76.480 ;
        RECT 71.960 76.410 72.190 76.480 ;
        RECT 71.575 76.335 72.190 76.410 ;
        RECT 73.895 76.335 74.125 76.480 ;
        RECT 75.095 76.335 75.325 76.480 ;
        RECT 70.320 76.165 75.325 76.335 ;
        RECT 70.320 76.020 70.550 76.165 ;
        RECT 71.575 76.090 72.190 76.165 ;
        RECT 71.960 76.020 72.190 76.090 ;
        RECT 73.895 76.020 74.125 76.165 ;
        RECT 75.095 76.020 75.325 76.165 ;
        RECT 75.530 76.135 75.820 77.210 ;
        RECT 70.755 75.880 71.755 75.910 ;
        RECT 74.285 75.880 74.935 75.910 ;
        RECT 75.525 75.880 75.825 76.135 ;
        RECT 70.735 75.710 71.775 75.880 ;
        RECT 74.265 75.775 75.825 75.880 ;
        RECT 74.265 75.710 75.820 75.775 ;
        RECT 70.755 75.680 71.755 75.710 ;
        RECT 74.285 75.680 74.935 75.710 ;
        RECT 71.170 75.320 71.340 75.680 ;
        RECT 70.755 75.290 71.755 75.320 ;
        RECT 72.890 75.290 73.150 75.365 ;
        RECT 74.285 75.290 74.935 75.320 ;
        RECT 70.735 75.120 71.775 75.290 ;
        RECT 72.890 75.120 74.955 75.290 ;
        RECT 70.755 75.090 71.755 75.120 ;
        RECT 72.890 75.045 73.150 75.120 ;
        RECT 74.285 75.090 74.935 75.120 ;
        RECT 70.320 74.835 70.550 74.980 ;
        RECT 71.960 74.910 72.190 74.980 ;
        RECT 71.960 74.835 72.255 74.910 ;
        RECT 73.895 74.835 74.125 74.980 ;
        RECT 75.095 74.835 75.325 74.980 ;
        RECT 70.320 74.665 75.325 74.835 ;
        RECT 63.155 74.275 65.065 74.380 ;
        RECT 50.625 72.880 51.625 72.910 ;
        RECT 54.155 72.880 54.805 72.910 ;
        RECT 55.395 72.880 55.695 73.135 ;
        RECT 50.605 72.710 51.645 72.880 ;
        RECT 54.135 72.775 55.695 72.880 ;
        RECT 54.135 72.710 55.690 72.775 ;
        RECT 50.625 72.680 51.625 72.710 ;
        RECT 54.155 72.680 54.805 72.710 ;
        RECT 51.040 72.320 51.210 72.680 ;
        RECT 50.625 72.290 51.625 72.320 ;
        RECT 52.760 72.290 53.020 72.365 ;
        RECT 54.155 72.290 54.805 72.320 ;
        RECT 50.605 72.120 51.645 72.290 ;
        RECT 52.760 72.120 54.825 72.290 ;
        RECT 50.625 72.090 51.625 72.120 ;
        RECT 52.760 72.045 53.020 72.120 ;
        RECT 54.155 72.090 54.805 72.120 ;
        RECT 50.190 71.835 50.420 71.980 ;
        RECT 51.025 71.835 51.285 71.910 ;
        RECT 51.830 71.835 52.060 71.980 ;
        RECT 53.765 71.835 53.995 71.980 ;
        RECT 54.965 71.835 55.195 71.980 ;
        RECT 50.190 71.665 55.195 71.835 ;
        RECT 37.205 71.180 38.205 71.210 ;
        RECT 40.735 71.180 41.385 71.210 ;
        RECT 37.620 70.820 37.790 71.180 ;
        RECT 37.205 70.790 38.205 70.820 ;
        RECT 39.340 70.790 39.600 70.865 ;
        RECT 40.735 70.790 41.385 70.820 ;
        RECT 37.185 70.620 38.225 70.790 ;
        RECT 39.340 70.620 41.405 70.790 ;
        RECT 37.205 70.590 38.205 70.620 ;
        RECT 39.340 70.545 39.600 70.620 ;
        RECT 40.735 70.590 41.385 70.620 ;
        RECT 36.770 70.335 37.000 70.480 ;
        RECT 38.410 70.410 38.640 70.480 ;
        RECT 38.410 70.335 38.705 70.410 ;
        RECT 40.345 70.335 40.575 70.480 ;
        RECT 41.545 70.335 41.775 70.480 ;
        RECT 36.770 70.165 41.775 70.335 ;
        RECT 36.770 70.020 37.000 70.165 ;
        RECT 38.410 70.090 38.705 70.165 ;
        RECT 38.410 70.020 38.640 70.090 ;
        RECT 40.345 70.020 40.575 70.165 ;
        RECT 41.545 70.020 41.775 70.165 ;
        RECT 41.980 70.135 42.270 71.210 ;
        RECT 37.205 69.880 38.205 69.910 ;
        RECT 40.735 69.880 41.385 69.910 ;
        RECT 41.975 69.880 42.275 70.135 ;
        RECT 36.320 69.710 38.225 69.880 ;
        RECT 40.715 69.775 42.275 69.880 ;
        RECT 43.030 69.880 43.320 71.275 ;
        RECT 43.895 71.210 44.935 71.380 ;
        RECT 47.425 71.210 48.980 71.380 ;
        RECT 49.735 71.275 50.035 71.635 ;
        RECT 50.190 71.520 50.420 71.665 ;
        RECT 51.025 71.590 51.285 71.665 ;
        RECT 51.830 71.520 52.060 71.665 ;
        RECT 53.765 71.520 53.995 71.665 ;
        RECT 54.965 71.520 55.195 71.665 ;
        RECT 50.625 71.380 51.625 71.410 ;
        RECT 54.155 71.380 54.805 71.410 ;
        RECT 55.400 71.380 55.690 72.710 ;
        RECT 56.450 71.635 56.740 74.210 ;
        RECT 57.335 74.180 58.335 74.210 ;
        RECT 60.865 74.180 61.515 74.210 ;
        RECT 57.335 73.790 58.335 73.820 ;
        RECT 59.470 73.790 59.730 73.865 ;
        RECT 60.865 73.790 61.515 73.820 ;
        RECT 57.315 73.620 61.535 73.790 ;
        RECT 57.335 73.590 58.335 73.620 ;
        RECT 59.470 73.545 59.730 73.620 ;
        RECT 60.865 73.590 61.515 73.620 ;
        RECT 56.900 73.335 57.130 73.480 ;
        RECT 57.315 73.335 57.575 73.410 ;
        RECT 58.540 73.335 58.770 73.480 ;
        RECT 60.475 73.335 60.705 73.480 ;
        RECT 61.675 73.335 61.905 73.480 ;
        RECT 56.900 73.165 61.905 73.335 ;
        RECT 56.900 73.020 57.130 73.165 ;
        RECT 57.315 73.090 57.575 73.165 ;
        RECT 58.540 73.020 58.770 73.165 ;
        RECT 60.475 73.020 60.705 73.165 ;
        RECT 61.675 73.020 61.905 73.165 ;
        RECT 62.110 73.135 62.400 74.210 ;
        RECT 63.160 74.210 65.065 74.275 ;
        RECT 67.555 74.210 69.110 74.380 ;
        RECT 69.865 74.380 70.165 74.635 ;
        RECT 70.320 74.520 70.550 74.665 ;
        RECT 71.960 74.590 72.255 74.665 ;
        RECT 71.960 74.520 72.190 74.590 ;
        RECT 73.895 74.520 74.125 74.665 ;
        RECT 75.095 74.520 75.325 74.665 ;
        RECT 70.755 74.380 71.755 74.410 ;
        RECT 74.285 74.380 74.935 74.410 ;
        RECT 75.530 74.380 75.820 75.710 ;
        RECT 76.580 74.635 76.870 77.275 ;
        RECT 77.445 77.210 78.485 77.380 ;
        RECT 80.975 77.210 82.530 77.380 ;
        RECT 83.285 77.275 83.585 77.635 ;
        RECT 83.740 77.520 83.970 77.665 ;
        RECT 84.155 77.590 84.415 77.665 ;
        RECT 85.380 77.520 85.610 77.665 ;
        RECT 87.315 77.520 87.545 77.665 ;
        RECT 88.515 77.520 88.745 77.665 ;
        RECT 84.175 77.380 85.175 77.410 ;
        RECT 87.705 77.380 88.355 77.410 ;
        RECT 88.950 77.380 89.240 78.500 ;
        RECT 90.000 77.635 90.290 78.500 ;
        RECT 90.885 78.290 91.885 78.320 ;
        RECT 93.020 78.290 93.280 78.365 ;
        RECT 94.415 78.290 95.065 78.320 ;
        RECT 90.865 78.120 95.085 78.290 ;
        RECT 90.885 78.090 91.885 78.120 ;
        RECT 93.020 78.045 93.280 78.120 ;
        RECT 94.415 78.090 95.065 78.120 ;
        RECT 90.450 77.835 90.680 77.980 ;
        RECT 90.865 77.835 91.125 77.910 ;
        RECT 92.090 77.835 92.320 77.980 ;
        RECT 94.025 77.835 94.255 77.980 ;
        RECT 95.225 77.835 95.455 77.980 ;
        RECT 90.450 77.665 95.455 77.835 ;
        RECT 77.465 77.180 78.465 77.210 ;
        RECT 80.995 77.180 81.645 77.210 ;
        RECT 77.880 76.820 78.050 77.180 ;
        RECT 77.465 76.790 78.465 76.820 ;
        RECT 79.600 76.790 79.860 76.865 ;
        RECT 80.995 76.790 81.645 76.820 ;
        RECT 77.445 76.620 78.485 76.790 ;
        RECT 79.600 76.620 81.665 76.790 ;
        RECT 77.465 76.590 78.465 76.620 ;
        RECT 79.600 76.545 79.860 76.620 ;
        RECT 80.995 76.590 81.645 76.620 ;
        RECT 77.030 76.335 77.260 76.480 ;
        RECT 78.670 76.410 78.900 76.480 ;
        RECT 78.285 76.335 78.900 76.410 ;
        RECT 80.605 76.335 80.835 76.480 ;
        RECT 81.805 76.335 82.035 76.480 ;
        RECT 77.030 76.165 82.035 76.335 ;
        RECT 77.030 76.020 77.260 76.165 ;
        RECT 78.285 76.090 78.900 76.165 ;
        RECT 78.670 76.020 78.900 76.090 ;
        RECT 80.605 76.020 80.835 76.165 ;
        RECT 81.805 76.020 82.035 76.165 ;
        RECT 82.240 76.135 82.530 77.210 ;
        RECT 77.465 75.880 78.465 75.910 ;
        RECT 80.995 75.880 81.645 75.910 ;
        RECT 82.235 75.880 82.535 76.135 ;
        RECT 77.445 75.710 78.485 75.880 ;
        RECT 80.975 75.775 82.535 75.880 ;
        RECT 80.975 75.710 82.530 75.775 ;
        RECT 77.465 75.680 78.465 75.710 ;
        RECT 80.995 75.680 81.645 75.710 ;
        RECT 77.880 75.320 78.050 75.680 ;
        RECT 77.465 75.290 78.465 75.320 ;
        RECT 79.600 75.290 79.860 75.365 ;
        RECT 80.995 75.290 81.645 75.320 ;
        RECT 77.445 75.120 78.485 75.290 ;
        RECT 79.600 75.120 81.665 75.290 ;
        RECT 77.465 75.090 78.465 75.120 ;
        RECT 79.600 75.045 79.860 75.120 ;
        RECT 80.995 75.090 81.645 75.120 ;
        RECT 77.030 74.835 77.260 74.980 ;
        RECT 78.670 74.910 78.900 74.980 ;
        RECT 78.670 74.835 78.965 74.910 ;
        RECT 80.605 74.835 80.835 74.980 ;
        RECT 81.805 74.835 82.035 74.980 ;
        RECT 77.030 74.665 82.035 74.835 ;
        RECT 69.865 74.275 71.775 74.380 ;
        RECT 57.335 72.880 58.335 72.910 ;
        RECT 60.865 72.880 61.515 72.910 ;
        RECT 62.105 72.880 62.405 73.135 ;
        RECT 57.315 72.710 58.355 72.880 ;
        RECT 60.845 72.775 62.405 72.880 ;
        RECT 60.845 72.710 62.400 72.775 ;
        RECT 57.335 72.680 58.335 72.710 ;
        RECT 60.865 72.680 61.515 72.710 ;
        RECT 57.750 72.320 57.920 72.680 ;
        RECT 57.335 72.290 58.335 72.320 ;
        RECT 59.470 72.290 59.730 72.365 ;
        RECT 60.865 72.290 61.515 72.320 ;
        RECT 57.315 72.120 58.355 72.290 ;
        RECT 59.470 72.120 61.535 72.290 ;
        RECT 57.335 72.090 58.335 72.120 ;
        RECT 59.470 72.045 59.730 72.120 ;
        RECT 60.865 72.090 61.515 72.120 ;
        RECT 56.900 71.835 57.130 71.980 ;
        RECT 57.735 71.835 57.995 71.910 ;
        RECT 58.540 71.835 58.770 71.980 ;
        RECT 60.475 71.835 60.705 71.980 ;
        RECT 61.675 71.835 61.905 71.980 ;
        RECT 56.900 71.665 61.905 71.835 ;
        RECT 43.915 71.180 44.915 71.210 ;
        RECT 47.445 71.180 48.095 71.210 ;
        RECT 44.330 70.820 44.500 71.180 ;
        RECT 43.915 70.790 44.915 70.820 ;
        RECT 46.050 70.790 46.310 70.865 ;
        RECT 47.445 70.790 48.095 70.820 ;
        RECT 43.895 70.620 44.935 70.790 ;
        RECT 46.050 70.620 48.115 70.790 ;
        RECT 43.915 70.590 44.915 70.620 ;
        RECT 46.050 70.545 46.310 70.620 ;
        RECT 47.445 70.590 48.095 70.620 ;
        RECT 43.480 70.335 43.710 70.480 ;
        RECT 45.120 70.410 45.350 70.480 ;
        RECT 45.120 70.335 45.415 70.410 ;
        RECT 47.055 70.335 47.285 70.480 ;
        RECT 48.255 70.335 48.485 70.480 ;
        RECT 43.480 70.165 48.485 70.335 ;
        RECT 43.480 70.020 43.710 70.165 ;
        RECT 45.120 70.090 45.415 70.165 ;
        RECT 45.120 70.020 45.350 70.090 ;
        RECT 47.055 70.020 47.285 70.165 ;
        RECT 48.255 70.020 48.485 70.165 ;
        RECT 48.690 70.135 48.980 71.210 ;
        RECT 43.915 69.880 44.915 69.910 ;
        RECT 47.445 69.880 48.095 69.910 ;
        RECT 48.685 69.880 48.985 70.135 ;
        RECT 40.715 69.710 42.270 69.775 ;
        RECT 36.320 68.635 36.610 69.710 ;
        RECT 37.205 69.680 38.205 69.710 ;
        RECT 40.735 69.680 41.385 69.710 ;
        RECT 41.145 69.320 41.405 69.365 ;
        RECT 37.205 69.290 38.205 69.320 ;
        RECT 40.735 69.290 41.405 69.320 ;
        RECT 37.185 69.120 41.405 69.290 ;
        RECT 37.205 69.090 38.205 69.120 ;
        RECT 40.735 69.090 41.405 69.120 ;
        RECT 41.145 69.045 41.405 69.090 ;
        RECT 36.770 68.835 37.000 68.980 ;
        RECT 38.410 68.835 38.640 68.980 ;
        RECT 39.340 68.835 39.600 68.910 ;
        RECT 40.345 68.835 40.575 68.980 ;
        RECT 41.545 68.835 41.775 68.980 ;
        RECT 36.770 68.665 41.775 68.835 ;
        RECT 36.315 68.380 36.615 68.635 ;
        RECT 36.770 68.520 37.000 68.665 ;
        RECT 38.410 68.520 38.640 68.665 ;
        RECT 39.340 68.590 39.600 68.665 ;
        RECT 40.345 68.520 40.575 68.665 ;
        RECT 41.545 68.520 41.775 68.665 ;
        RECT 37.205 68.380 38.205 68.410 ;
        RECT 40.735 68.380 41.385 68.410 ;
        RECT 41.980 68.380 42.270 69.710 ;
        RECT 43.030 69.710 44.935 69.880 ;
        RECT 47.425 69.775 48.985 69.880 ;
        RECT 49.740 69.880 50.030 71.275 ;
        RECT 50.605 71.210 51.645 71.380 ;
        RECT 54.135 71.210 55.690 71.380 ;
        RECT 56.445 71.275 56.745 71.635 ;
        RECT 56.900 71.520 57.130 71.665 ;
        RECT 57.735 71.590 57.995 71.665 ;
        RECT 58.540 71.520 58.770 71.665 ;
        RECT 60.475 71.520 60.705 71.665 ;
        RECT 61.675 71.520 61.905 71.665 ;
        RECT 57.335 71.380 58.335 71.410 ;
        RECT 60.865 71.380 61.515 71.410 ;
        RECT 62.110 71.380 62.400 72.710 ;
        RECT 63.160 71.635 63.450 74.210 ;
        RECT 64.045 74.180 65.045 74.210 ;
        RECT 67.575 74.180 68.225 74.210 ;
        RECT 64.045 73.790 65.045 73.820 ;
        RECT 66.180 73.790 66.440 73.865 ;
        RECT 67.575 73.790 68.225 73.820 ;
        RECT 64.025 73.620 68.245 73.790 ;
        RECT 64.045 73.590 65.045 73.620 ;
        RECT 66.180 73.545 66.440 73.620 ;
        RECT 67.575 73.590 68.225 73.620 ;
        RECT 63.610 73.335 63.840 73.480 ;
        RECT 64.025 73.335 64.285 73.410 ;
        RECT 65.250 73.335 65.480 73.480 ;
        RECT 67.185 73.335 67.415 73.480 ;
        RECT 68.385 73.335 68.615 73.480 ;
        RECT 63.610 73.165 68.615 73.335 ;
        RECT 63.610 73.020 63.840 73.165 ;
        RECT 64.025 73.090 64.285 73.165 ;
        RECT 65.250 73.020 65.480 73.165 ;
        RECT 67.185 73.020 67.415 73.165 ;
        RECT 68.385 73.020 68.615 73.165 ;
        RECT 68.820 73.135 69.110 74.210 ;
        RECT 69.870 74.210 71.775 74.275 ;
        RECT 74.265 74.210 75.820 74.380 ;
        RECT 76.575 74.380 76.875 74.635 ;
        RECT 77.030 74.520 77.260 74.665 ;
        RECT 78.670 74.590 78.965 74.665 ;
        RECT 78.670 74.520 78.900 74.590 ;
        RECT 80.605 74.520 80.835 74.665 ;
        RECT 81.805 74.520 82.035 74.665 ;
        RECT 77.465 74.380 78.465 74.410 ;
        RECT 80.995 74.380 81.645 74.410 ;
        RECT 82.240 74.380 82.530 75.710 ;
        RECT 83.290 74.635 83.580 77.275 ;
        RECT 84.155 77.210 85.195 77.380 ;
        RECT 87.685 77.210 89.240 77.380 ;
        RECT 89.995 77.275 90.295 77.635 ;
        RECT 90.450 77.520 90.680 77.665 ;
        RECT 90.865 77.590 91.125 77.665 ;
        RECT 92.090 77.520 92.320 77.665 ;
        RECT 94.025 77.520 94.255 77.665 ;
        RECT 95.225 77.520 95.455 77.665 ;
        RECT 90.885 77.380 91.885 77.410 ;
        RECT 94.415 77.380 95.065 77.410 ;
        RECT 95.660 77.380 95.950 78.500 ;
        RECT 96.710 77.635 97.000 78.500 ;
        RECT 97.595 78.290 98.595 78.320 ;
        RECT 99.730 78.290 99.990 78.365 ;
        RECT 101.125 78.290 101.775 78.320 ;
        RECT 97.575 78.120 101.795 78.290 ;
        RECT 97.595 78.090 98.595 78.120 ;
        RECT 99.730 78.045 99.990 78.120 ;
        RECT 101.125 78.090 101.775 78.120 ;
        RECT 97.160 77.835 97.390 77.980 ;
        RECT 97.575 77.835 97.835 77.910 ;
        RECT 98.800 77.835 99.030 77.980 ;
        RECT 100.735 77.835 100.965 77.980 ;
        RECT 101.935 77.835 102.165 77.980 ;
        RECT 97.160 77.665 102.165 77.835 ;
        RECT 84.175 77.180 85.175 77.210 ;
        RECT 87.705 77.180 88.355 77.210 ;
        RECT 84.590 76.820 84.760 77.180 ;
        RECT 84.175 76.790 85.175 76.820 ;
        RECT 86.310 76.790 86.570 76.865 ;
        RECT 87.705 76.790 88.355 76.820 ;
        RECT 84.155 76.620 85.195 76.790 ;
        RECT 86.310 76.620 88.375 76.790 ;
        RECT 84.175 76.590 85.175 76.620 ;
        RECT 86.310 76.545 86.570 76.620 ;
        RECT 87.705 76.590 88.355 76.620 ;
        RECT 83.740 76.335 83.970 76.480 ;
        RECT 85.380 76.410 85.610 76.480 ;
        RECT 84.995 76.335 85.610 76.410 ;
        RECT 87.315 76.335 87.545 76.480 ;
        RECT 88.515 76.335 88.745 76.480 ;
        RECT 83.740 76.165 88.745 76.335 ;
        RECT 83.740 76.020 83.970 76.165 ;
        RECT 84.995 76.090 85.610 76.165 ;
        RECT 85.380 76.020 85.610 76.090 ;
        RECT 87.315 76.020 87.545 76.165 ;
        RECT 88.515 76.020 88.745 76.165 ;
        RECT 88.950 76.135 89.240 77.210 ;
        RECT 84.175 75.880 85.175 75.910 ;
        RECT 87.705 75.880 88.355 75.910 ;
        RECT 88.945 75.880 89.245 76.135 ;
        RECT 84.155 75.710 85.195 75.880 ;
        RECT 87.685 75.775 89.245 75.880 ;
        RECT 87.685 75.710 89.240 75.775 ;
        RECT 84.175 75.680 85.175 75.710 ;
        RECT 87.705 75.680 88.355 75.710 ;
        RECT 84.590 75.320 84.760 75.680 ;
        RECT 84.175 75.290 85.175 75.320 ;
        RECT 86.310 75.290 86.570 75.365 ;
        RECT 87.705 75.290 88.355 75.320 ;
        RECT 84.155 75.120 85.195 75.290 ;
        RECT 86.310 75.120 88.375 75.290 ;
        RECT 84.175 75.090 85.175 75.120 ;
        RECT 86.310 75.045 86.570 75.120 ;
        RECT 87.705 75.090 88.355 75.120 ;
        RECT 83.740 74.835 83.970 74.980 ;
        RECT 85.380 74.910 85.610 74.980 ;
        RECT 85.380 74.835 85.675 74.910 ;
        RECT 87.315 74.835 87.545 74.980 ;
        RECT 88.515 74.835 88.745 74.980 ;
        RECT 83.740 74.665 88.745 74.835 ;
        RECT 76.575 74.275 78.485 74.380 ;
        RECT 64.045 72.880 65.045 72.910 ;
        RECT 67.575 72.880 68.225 72.910 ;
        RECT 68.815 72.880 69.115 73.135 ;
        RECT 64.025 72.710 65.065 72.880 ;
        RECT 67.555 72.775 69.115 72.880 ;
        RECT 67.555 72.710 69.110 72.775 ;
        RECT 64.045 72.680 65.045 72.710 ;
        RECT 67.575 72.680 68.225 72.710 ;
        RECT 64.460 72.320 64.630 72.680 ;
        RECT 64.045 72.290 65.045 72.320 ;
        RECT 66.180 72.290 66.440 72.365 ;
        RECT 67.575 72.290 68.225 72.320 ;
        RECT 64.025 72.120 65.065 72.290 ;
        RECT 66.180 72.120 68.245 72.290 ;
        RECT 64.045 72.090 65.045 72.120 ;
        RECT 66.180 72.045 66.440 72.120 ;
        RECT 67.575 72.090 68.225 72.120 ;
        RECT 63.610 71.835 63.840 71.980 ;
        RECT 64.445 71.835 64.705 71.910 ;
        RECT 65.250 71.835 65.480 71.980 ;
        RECT 67.185 71.835 67.415 71.980 ;
        RECT 68.385 71.835 68.615 71.980 ;
        RECT 63.610 71.665 68.615 71.835 ;
        RECT 50.625 71.180 51.625 71.210 ;
        RECT 54.155 71.180 54.805 71.210 ;
        RECT 51.040 70.820 51.210 71.180 ;
        RECT 50.625 70.790 51.625 70.820 ;
        RECT 52.760 70.790 53.020 70.865 ;
        RECT 54.155 70.790 54.805 70.820 ;
        RECT 50.605 70.620 51.645 70.790 ;
        RECT 52.760 70.620 54.825 70.790 ;
        RECT 50.625 70.590 51.625 70.620 ;
        RECT 52.760 70.545 53.020 70.620 ;
        RECT 54.155 70.590 54.805 70.620 ;
        RECT 50.190 70.335 50.420 70.480 ;
        RECT 51.830 70.410 52.060 70.480 ;
        RECT 51.830 70.335 52.125 70.410 ;
        RECT 53.765 70.335 53.995 70.480 ;
        RECT 54.965 70.335 55.195 70.480 ;
        RECT 50.190 70.165 55.195 70.335 ;
        RECT 50.190 70.020 50.420 70.165 ;
        RECT 51.830 70.090 52.125 70.165 ;
        RECT 51.830 70.020 52.060 70.090 ;
        RECT 53.765 70.020 53.995 70.165 ;
        RECT 54.965 70.020 55.195 70.165 ;
        RECT 55.400 70.135 55.690 71.210 ;
        RECT 50.625 69.880 51.625 69.910 ;
        RECT 54.155 69.880 54.805 69.910 ;
        RECT 55.395 69.880 55.695 70.135 ;
        RECT 47.425 69.710 48.980 69.775 ;
        RECT 43.030 68.635 43.320 69.710 ;
        RECT 43.915 69.680 44.915 69.710 ;
        RECT 47.445 69.680 48.095 69.710 ;
        RECT 44.315 69.320 44.575 69.365 ;
        RECT 43.915 69.290 44.915 69.320 ;
        RECT 47.445 69.290 48.095 69.320 ;
        RECT 43.895 69.120 48.115 69.290 ;
        RECT 43.915 69.090 44.915 69.120 ;
        RECT 47.445 69.090 48.095 69.120 ;
        RECT 44.315 69.045 44.575 69.090 ;
        RECT 43.480 68.835 43.710 68.980 ;
        RECT 45.120 68.835 45.350 68.980 ;
        RECT 46.050 68.835 46.310 68.910 ;
        RECT 47.055 68.835 47.285 68.980 ;
        RECT 48.255 68.835 48.485 68.980 ;
        RECT 43.480 68.665 48.485 68.835 ;
        RECT 36.315 68.275 38.225 68.380 ;
        RECT 36.320 68.210 38.225 68.275 ;
        RECT 36.320 66.880 36.610 68.210 ;
        RECT 37.205 68.180 38.205 68.210 ;
        RECT 38.450 67.950 38.710 68.270 ;
        RECT 40.715 68.210 42.270 68.380 ;
        RECT 43.025 68.380 43.325 68.635 ;
        RECT 43.480 68.520 43.710 68.665 ;
        RECT 45.120 68.520 45.350 68.665 ;
        RECT 46.050 68.590 46.310 68.665 ;
        RECT 47.055 68.520 47.285 68.665 ;
        RECT 48.255 68.520 48.485 68.665 ;
        RECT 43.915 68.380 44.915 68.410 ;
        RECT 47.445 68.380 48.095 68.410 ;
        RECT 48.690 68.380 48.980 69.710 ;
        RECT 49.740 69.710 51.645 69.880 ;
        RECT 54.135 69.775 55.695 69.880 ;
        RECT 56.450 69.880 56.740 71.275 ;
        RECT 57.315 71.210 58.355 71.380 ;
        RECT 60.845 71.210 62.400 71.380 ;
        RECT 63.155 71.275 63.455 71.635 ;
        RECT 63.610 71.520 63.840 71.665 ;
        RECT 64.445 71.590 64.705 71.665 ;
        RECT 65.250 71.520 65.480 71.665 ;
        RECT 67.185 71.520 67.415 71.665 ;
        RECT 68.385 71.520 68.615 71.665 ;
        RECT 64.045 71.380 65.045 71.410 ;
        RECT 67.575 71.380 68.225 71.410 ;
        RECT 68.820 71.380 69.110 72.710 ;
        RECT 69.870 71.635 70.160 74.210 ;
        RECT 70.755 74.180 71.755 74.210 ;
        RECT 74.285 74.180 74.935 74.210 ;
        RECT 70.755 73.790 71.755 73.820 ;
        RECT 72.890 73.790 73.150 73.865 ;
        RECT 74.285 73.790 74.935 73.820 ;
        RECT 70.735 73.620 74.955 73.790 ;
        RECT 70.755 73.590 71.755 73.620 ;
        RECT 72.890 73.545 73.150 73.620 ;
        RECT 74.285 73.590 74.935 73.620 ;
        RECT 70.320 73.335 70.550 73.480 ;
        RECT 70.735 73.335 70.995 73.410 ;
        RECT 71.960 73.335 72.190 73.480 ;
        RECT 73.895 73.335 74.125 73.480 ;
        RECT 75.095 73.335 75.325 73.480 ;
        RECT 70.320 73.165 75.325 73.335 ;
        RECT 70.320 73.020 70.550 73.165 ;
        RECT 70.735 73.090 70.995 73.165 ;
        RECT 71.960 73.020 72.190 73.165 ;
        RECT 73.895 73.020 74.125 73.165 ;
        RECT 75.095 73.020 75.325 73.165 ;
        RECT 75.530 73.135 75.820 74.210 ;
        RECT 76.580 74.210 78.485 74.275 ;
        RECT 80.975 74.210 82.530 74.380 ;
        RECT 83.285 74.380 83.585 74.635 ;
        RECT 83.740 74.520 83.970 74.665 ;
        RECT 85.380 74.590 85.675 74.665 ;
        RECT 85.380 74.520 85.610 74.590 ;
        RECT 87.315 74.520 87.545 74.665 ;
        RECT 88.515 74.520 88.745 74.665 ;
        RECT 84.175 74.380 85.175 74.410 ;
        RECT 87.705 74.380 88.355 74.410 ;
        RECT 88.950 74.380 89.240 75.710 ;
        RECT 90.000 74.635 90.290 77.275 ;
        RECT 90.865 77.210 91.905 77.380 ;
        RECT 94.395 77.210 95.950 77.380 ;
        RECT 96.705 77.275 97.005 77.635 ;
        RECT 97.160 77.520 97.390 77.665 ;
        RECT 97.575 77.590 97.835 77.665 ;
        RECT 98.800 77.520 99.030 77.665 ;
        RECT 100.735 77.520 100.965 77.665 ;
        RECT 101.935 77.520 102.165 77.665 ;
        RECT 97.595 77.380 98.595 77.410 ;
        RECT 101.125 77.380 101.775 77.410 ;
        RECT 102.370 77.380 102.660 78.500 ;
        RECT 90.885 77.180 91.885 77.210 ;
        RECT 94.415 77.180 95.065 77.210 ;
        RECT 91.300 76.820 91.470 77.180 ;
        RECT 90.885 76.790 91.885 76.820 ;
        RECT 93.020 76.790 93.280 76.865 ;
        RECT 94.415 76.790 95.065 76.820 ;
        RECT 90.865 76.620 91.905 76.790 ;
        RECT 93.020 76.620 95.085 76.790 ;
        RECT 90.885 76.590 91.885 76.620 ;
        RECT 93.020 76.545 93.280 76.620 ;
        RECT 94.415 76.590 95.065 76.620 ;
        RECT 90.450 76.335 90.680 76.480 ;
        RECT 92.090 76.410 92.320 76.480 ;
        RECT 91.705 76.335 92.320 76.410 ;
        RECT 94.025 76.335 94.255 76.480 ;
        RECT 95.225 76.335 95.455 76.480 ;
        RECT 90.450 76.165 95.455 76.335 ;
        RECT 90.450 76.020 90.680 76.165 ;
        RECT 91.705 76.090 92.320 76.165 ;
        RECT 92.090 76.020 92.320 76.090 ;
        RECT 94.025 76.020 94.255 76.165 ;
        RECT 95.225 76.020 95.455 76.165 ;
        RECT 95.660 76.135 95.950 77.210 ;
        RECT 90.885 75.880 91.885 75.910 ;
        RECT 94.415 75.880 95.065 75.910 ;
        RECT 95.655 75.880 95.955 76.135 ;
        RECT 90.865 75.710 91.905 75.880 ;
        RECT 94.395 75.775 95.955 75.880 ;
        RECT 94.395 75.710 95.950 75.775 ;
        RECT 90.885 75.680 91.885 75.710 ;
        RECT 94.415 75.680 95.065 75.710 ;
        RECT 91.300 75.320 91.470 75.680 ;
        RECT 90.885 75.290 91.885 75.320 ;
        RECT 93.020 75.290 93.280 75.365 ;
        RECT 94.415 75.290 95.065 75.320 ;
        RECT 90.865 75.120 91.905 75.290 ;
        RECT 93.020 75.120 95.085 75.290 ;
        RECT 90.885 75.090 91.885 75.120 ;
        RECT 93.020 75.045 93.280 75.120 ;
        RECT 94.415 75.090 95.065 75.120 ;
        RECT 90.450 74.835 90.680 74.980 ;
        RECT 92.090 74.910 92.320 74.980 ;
        RECT 92.090 74.835 92.385 74.910 ;
        RECT 94.025 74.835 94.255 74.980 ;
        RECT 95.225 74.835 95.455 74.980 ;
        RECT 90.450 74.665 95.455 74.835 ;
        RECT 83.285 74.275 85.195 74.380 ;
        RECT 70.755 72.880 71.755 72.910 ;
        RECT 74.285 72.880 74.935 72.910 ;
        RECT 75.525 72.880 75.825 73.135 ;
        RECT 70.735 72.710 71.775 72.880 ;
        RECT 74.265 72.775 75.825 72.880 ;
        RECT 74.265 72.710 75.820 72.775 ;
        RECT 70.755 72.680 71.755 72.710 ;
        RECT 74.285 72.680 74.935 72.710 ;
        RECT 71.170 72.320 71.340 72.680 ;
        RECT 70.755 72.290 71.755 72.320 ;
        RECT 72.890 72.290 73.150 72.365 ;
        RECT 74.285 72.290 74.935 72.320 ;
        RECT 70.735 72.120 71.775 72.290 ;
        RECT 72.890 72.120 74.955 72.290 ;
        RECT 70.755 72.090 71.755 72.120 ;
        RECT 72.890 72.045 73.150 72.120 ;
        RECT 74.285 72.090 74.935 72.120 ;
        RECT 70.320 71.835 70.550 71.980 ;
        RECT 71.155 71.835 71.415 71.910 ;
        RECT 71.960 71.835 72.190 71.980 ;
        RECT 73.895 71.835 74.125 71.980 ;
        RECT 75.095 71.835 75.325 71.980 ;
        RECT 70.320 71.665 75.325 71.835 ;
        RECT 57.335 71.180 58.335 71.210 ;
        RECT 60.865 71.180 61.515 71.210 ;
        RECT 57.750 70.820 57.920 71.180 ;
        RECT 57.335 70.790 58.335 70.820 ;
        RECT 59.470 70.790 59.730 70.865 ;
        RECT 60.865 70.790 61.515 70.820 ;
        RECT 57.315 70.620 58.355 70.790 ;
        RECT 59.470 70.620 61.535 70.790 ;
        RECT 57.335 70.590 58.335 70.620 ;
        RECT 59.470 70.545 59.730 70.620 ;
        RECT 60.865 70.590 61.515 70.620 ;
        RECT 56.900 70.335 57.130 70.480 ;
        RECT 58.540 70.410 58.770 70.480 ;
        RECT 58.540 70.335 58.835 70.410 ;
        RECT 60.475 70.335 60.705 70.480 ;
        RECT 61.675 70.335 61.905 70.480 ;
        RECT 56.900 70.165 61.905 70.335 ;
        RECT 56.900 70.020 57.130 70.165 ;
        RECT 58.540 70.090 58.835 70.165 ;
        RECT 58.540 70.020 58.770 70.090 ;
        RECT 60.475 70.020 60.705 70.165 ;
        RECT 61.675 70.020 61.905 70.165 ;
        RECT 62.110 70.135 62.400 71.210 ;
        RECT 57.335 69.880 58.335 69.910 ;
        RECT 60.865 69.880 61.515 69.910 ;
        RECT 62.105 69.880 62.405 70.135 ;
        RECT 54.135 69.710 55.690 69.775 ;
        RECT 49.740 68.635 50.030 69.710 ;
        RECT 50.625 69.680 51.625 69.710 ;
        RECT 54.155 69.680 54.805 69.710 ;
        RECT 54.565 69.320 54.825 69.365 ;
        RECT 50.625 69.290 51.625 69.320 ;
        RECT 54.155 69.290 54.825 69.320 ;
        RECT 50.605 69.120 54.825 69.290 ;
        RECT 50.625 69.090 51.625 69.120 ;
        RECT 54.155 69.090 54.825 69.120 ;
        RECT 54.565 69.045 54.825 69.090 ;
        RECT 50.190 68.835 50.420 68.980 ;
        RECT 51.830 68.835 52.060 68.980 ;
        RECT 52.760 68.835 53.020 68.910 ;
        RECT 53.765 68.835 53.995 68.980 ;
        RECT 54.965 68.835 55.195 68.980 ;
        RECT 50.190 68.665 55.195 68.835 ;
        RECT 43.025 68.275 44.935 68.380 ;
        RECT 40.735 68.180 41.385 68.210 ;
        RECT 37.205 67.790 38.205 67.820 ;
        RECT 38.495 67.790 38.665 67.950 ;
        RECT 39.340 67.790 39.600 67.865 ;
        RECT 40.735 67.790 41.385 67.820 ;
        RECT 37.185 67.620 41.405 67.790 ;
        RECT 37.205 67.590 38.205 67.620 ;
        RECT 39.340 67.545 39.600 67.620 ;
        RECT 40.735 67.590 41.385 67.620 ;
        RECT 36.770 67.335 37.000 67.480 ;
        RECT 38.410 67.335 38.640 67.480 ;
        RECT 39.310 67.335 39.630 67.380 ;
        RECT 40.345 67.335 40.575 67.480 ;
        RECT 41.545 67.335 41.775 67.480 ;
        RECT 36.770 67.165 41.775 67.335 ;
        RECT 36.770 67.020 37.000 67.165 ;
        RECT 38.410 67.020 38.640 67.165 ;
        RECT 39.310 67.120 39.630 67.165 ;
        RECT 40.345 67.020 40.575 67.165 ;
        RECT 41.545 67.020 41.775 67.165 ;
        RECT 41.980 67.135 42.270 68.210 ;
        RECT 43.030 68.210 44.935 68.275 ;
        RECT 47.425 68.210 48.980 68.380 ;
        RECT 49.735 68.380 50.035 68.635 ;
        RECT 50.190 68.520 50.420 68.665 ;
        RECT 51.830 68.520 52.060 68.665 ;
        RECT 52.760 68.590 53.020 68.665 ;
        RECT 53.765 68.520 53.995 68.665 ;
        RECT 54.965 68.520 55.195 68.665 ;
        RECT 50.625 68.380 51.625 68.410 ;
        RECT 54.155 68.380 54.805 68.410 ;
        RECT 55.400 68.380 55.690 69.710 ;
        RECT 56.450 69.710 58.355 69.880 ;
        RECT 60.845 69.775 62.405 69.880 ;
        RECT 63.160 69.880 63.450 71.275 ;
        RECT 64.025 71.210 65.065 71.380 ;
        RECT 67.555 71.210 69.110 71.380 ;
        RECT 69.865 71.275 70.165 71.635 ;
        RECT 70.320 71.520 70.550 71.665 ;
        RECT 71.155 71.590 71.415 71.665 ;
        RECT 71.960 71.520 72.190 71.665 ;
        RECT 73.895 71.520 74.125 71.665 ;
        RECT 75.095 71.520 75.325 71.665 ;
        RECT 70.755 71.380 71.755 71.410 ;
        RECT 74.285 71.380 74.935 71.410 ;
        RECT 75.530 71.380 75.820 72.710 ;
        RECT 76.580 71.635 76.870 74.210 ;
        RECT 77.465 74.180 78.465 74.210 ;
        RECT 80.995 74.180 81.645 74.210 ;
        RECT 77.465 73.790 78.465 73.820 ;
        RECT 79.600 73.790 79.860 73.865 ;
        RECT 80.995 73.790 81.645 73.820 ;
        RECT 77.445 73.620 81.665 73.790 ;
        RECT 77.465 73.590 78.465 73.620 ;
        RECT 79.600 73.545 79.860 73.620 ;
        RECT 80.995 73.590 81.645 73.620 ;
        RECT 77.030 73.335 77.260 73.480 ;
        RECT 77.445 73.335 77.705 73.410 ;
        RECT 78.670 73.335 78.900 73.480 ;
        RECT 80.605 73.335 80.835 73.480 ;
        RECT 81.805 73.335 82.035 73.480 ;
        RECT 77.030 73.165 82.035 73.335 ;
        RECT 77.030 73.020 77.260 73.165 ;
        RECT 77.445 73.090 77.705 73.165 ;
        RECT 78.670 73.020 78.900 73.165 ;
        RECT 80.605 73.020 80.835 73.165 ;
        RECT 81.805 73.020 82.035 73.165 ;
        RECT 82.240 73.135 82.530 74.210 ;
        RECT 83.290 74.210 85.195 74.275 ;
        RECT 87.685 74.210 89.240 74.380 ;
        RECT 89.995 74.380 90.295 74.635 ;
        RECT 90.450 74.520 90.680 74.665 ;
        RECT 92.090 74.590 92.385 74.665 ;
        RECT 92.090 74.520 92.320 74.590 ;
        RECT 94.025 74.520 94.255 74.665 ;
        RECT 95.225 74.520 95.455 74.665 ;
        RECT 90.885 74.380 91.885 74.410 ;
        RECT 94.415 74.380 95.065 74.410 ;
        RECT 95.660 74.380 95.950 75.710 ;
        RECT 96.710 74.635 97.000 77.275 ;
        RECT 97.575 77.210 98.615 77.380 ;
        RECT 101.105 77.210 102.660 77.380 ;
        RECT 97.595 77.180 98.595 77.210 ;
        RECT 101.125 77.180 101.775 77.210 ;
        RECT 98.010 76.820 98.180 77.180 ;
        RECT 97.595 76.790 98.595 76.820 ;
        RECT 99.730 76.790 99.990 76.865 ;
        RECT 101.125 76.790 101.775 76.820 ;
        RECT 97.575 76.620 98.615 76.790 ;
        RECT 99.730 76.620 101.795 76.790 ;
        RECT 97.595 76.590 98.595 76.620 ;
        RECT 99.730 76.545 99.990 76.620 ;
        RECT 101.125 76.590 101.775 76.620 ;
        RECT 97.160 76.335 97.390 76.480 ;
        RECT 98.800 76.410 99.030 76.480 ;
        RECT 98.415 76.335 99.030 76.410 ;
        RECT 100.735 76.335 100.965 76.480 ;
        RECT 101.935 76.335 102.165 76.480 ;
        RECT 97.160 76.165 102.165 76.335 ;
        RECT 97.160 76.020 97.390 76.165 ;
        RECT 98.415 76.090 99.030 76.165 ;
        RECT 98.800 76.020 99.030 76.090 ;
        RECT 100.735 76.020 100.965 76.165 ;
        RECT 101.935 76.020 102.165 76.165 ;
        RECT 102.370 76.135 102.660 77.210 ;
        RECT 97.595 75.880 98.595 75.910 ;
        RECT 101.125 75.880 101.775 75.910 ;
        RECT 102.365 75.880 102.665 76.135 ;
        RECT 97.575 75.710 98.615 75.880 ;
        RECT 101.105 75.775 102.665 75.880 ;
        RECT 101.105 75.710 102.660 75.775 ;
        RECT 97.595 75.680 98.595 75.710 ;
        RECT 101.125 75.680 101.775 75.710 ;
        RECT 98.010 75.320 98.180 75.680 ;
        RECT 97.595 75.290 98.595 75.320 ;
        RECT 99.730 75.290 99.990 75.365 ;
        RECT 101.125 75.290 101.775 75.320 ;
        RECT 97.575 75.120 98.615 75.290 ;
        RECT 99.730 75.120 101.795 75.290 ;
        RECT 97.595 75.090 98.595 75.120 ;
        RECT 99.730 75.045 99.990 75.120 ;
        RECT 101.125 75.090 101.775 75.120 ;
        RECT 97.160 74.835 97.390 74.980 ;
        RECT 98.800 74.910 99.030 74.980 ;
        RECT 98.800 74.835 99.095 74.910 ;
        RECT 100.735 74.835 100.965 74.980 ;
        RECT 101.935 74.835 102.165 74.980 ;
        RECT 97.160 74.665 102.165 74.835 ;
        RECT 89.995 74.275 91.905 74.380 ;
        RECT 77.465 72.880 78.465 72.910 ;
        RECT 80.995 72.880 81.645 72.910 ;
        RECT 82.235 72.880 82.535 73.135 ;
        RECT 77.445 72.710 78.485 72.880 ;
        RECT 80.975 72.775 82.535 72.880 ;
        RECT 80.975 72.710 82.530 72.775 ;
        RECT 77.465 72.680 78.465 72.710 ;
        RECT 80.995 72.680 81.645 72.710 ;
        RECT 77.880 72.320 78.050 72.680 ;
        RECT 77.465 72.290 78.465 72.320 ;
        RECT 79.600 72.290 79.860 72.365 ;
        RECT 80.995 72.290 81.645 72.320 ;
        RECT 77.445 72.120 78.485 72.290 ;
        RECT 79.600 72.120 81.665 72.290 ;
        RECT 77.465 72.090 78.465 72.120 ;
        RECT 79.600 72.045 79.860 72.120 ;
        RECT 80.995 72.090 81.645 72.120 ;
        RECT 77.030 71.835 77.260 71.980 ;
        RECT 77.865 71.835 78.125 71.910 ;
        RECT 78.670 71.835 78.900 71.980 ;
        RECT 80.605 71.835 80.835 71.980 ;
        RECT 81.805 71.835 82.035 71.980 ;
        RECT 77.030 71.665 82.035 71.835 ;
        RECT 64.045 71.180 65.045 71.210 ;
        RECT 67.575 71.180 68.225 71.210 ;
        RECT 64.460 70.820 64.630 71.180 ;
        RECT 64.045 70.790 65.045 70.820 ;
        RECT 66.180 70.790 66.440 70.865 ;
        RECT 67.575 70.790 68.225 70.820 ;
        RECT 64.025 70.620 65.065 70.790 ;
        RECT 66.180 70.620 68.245 70.790 ;
        RECT 64.045 70.590 65.045 70.620 ;
        RECT 66.180 70.545 66.440 70.620 ;
        RECT 67.575 70.590 68.225 70.620 ;
        RECT 63.610 70.335 63.840 70.480 ;
        RECT 65.250 70.410 65.480 70.480 ;
        RECT 65.250 70.335 65.545 70.410 ;
        RECT 67.185 70.335 67.415 70.480 ;
        RECT 68.385 70.335 68.615 70.480 ;
        RECT 63.610 70.165 68.615 70.335 ;
        RECT 63.610 70.020 63.840 70.165 ;
        RECT 65.250 70.090 65.545 70.165 ;
        RECT 65.250 70.020 65.480 70.090 ;
        RECT 67.185 70.020 67.415 70.165 ;
        RECT 68.385 70.020 68.615 70.165 ;
        RECT 68.820 70.135 69.110 71.210 ;
        RECT 64.045 69.880 65.045 69.910 ;
        RECT 67.575 69.880 68.225 69.910 ;
        RECT 68.815 69.880 69.115 70.135 ;
        RECT 60.845 69.710 62.400 69.775 ;
        RECT 56.450 68.635 56.740 69.710 ;
        RECT 57.335 69.680 58.335 69.710 ;
        RECT 60.865 69.680 61.515 69.710 ;
        RECT 57.735 69.320 57.995 69.365 ;
        RECT 57.335 69.290 58.335 69.320 ;
        RECT 60.865 69.290 61.515 69.320 ;
        RECT 57.315 69.120 61.535 69.290 ;
        RECT 57.335 69.090 58.335 69.120 ;
        RECT 60.865 69.090 61.515 69.120 ;
        RECT 57.735 69.045 57.995 69.090 ;
        RECT 56.900 68.835 57.130 68.980 ;
        RECT 58.540 68.835 58.770 68.980 ;
        RECT 59.470 68.835 59.730 68.910 ;
        RECT 60.475 68.835 60.705 68.980 ;
        RECT 61.675 68.835 61.905 68.980 ;
        RECT 56.900 68.665 61.905 68.835 ;
        RECT 49.735 68.275 51.645 68.380 ;
        RECT 37.205 66.880 38.205 66.910 ;
        RECT 40.735 66.880 41.385 66.910 ;
        RECT 41.975 66.880 42.275 67.135 ;
        RECT 36.320 66.710 38.225 66.880 ;
        RECT 40.715 66.775 42.275 66.880 ;
        RECT 43.030 66.880 43.320 68.210 ;
        RECT 43.915 68.180 44.915 68.210 ;
        RECT 47.445 68.180 48.095 68.210 ;
        RECT 44.735 67.820 44.995 67.865 ;
        RECT 43.915 67.790 44.995 67.820 ;
        RECT 46.050 67.790 46.310 67.865 ;
        RECT 47.445 67.790 48.095 67.820 ;
        RECT 43.895 67.620 48.115 67.790 ;
        RECT 43.915 67.590 44.995 67.620 ;
        RECT 44.735 67.545 44.995 67.590 ;
        RECT 46.050 67.545 46.310 67.620 ;
        RECT 47.445 67.590 48.095 67.620 ;
        RECT 43.480 67.335 43.710 67.480 ;
        RECT 45.120 67.335 45.350 67.480 ;
        RECT 46.020 67.335 46.340 67.380 ;
        RECT 47.055 67.335 47.285 67.480 ;
        RECT 48.255 67.335 48.485 67.480 ;
        RECT 43.480 67.165 48.485 67.335 ;
        RECT 43.480 67.020 43.710 67.165 ;
        RECT 45.120 67.020 45.350 67.165 ;
        RECT 46.020 67.120 46.340 67.165 ;
        RECT 47.055 67.020 47.285 67.165 ;
        RECT 48.255 67.020 48.485 67.165 ;
        RECT 48.690 67.135 48.980 68.210 ;
        RECT 49.740 68.210 51.645 68.275 ;
        RECT 43.915 66.880 44.915 66.910 ;
        RECT 47.445 66.880 48.095 66.910 ;
        RECT 48.685 66.880 48.985 67.135 ;
        RECT 40.715 66.710 42.270 66.775 ;
        RECT 36.320 65.635 36.610 66.710 ;
        RECT 37.205 66.680 38.205 66.710 ;
        RECT 40.735 66.680 41.385 66.710 ;
        RECT 37.205 66.290 38.205 66.320 ;
        RECT 40.735 66.290 41.385 66.320 ;
        RECT 37.185 66.120 41.405 66.290 ;
        RECT 37.205 66.090 38.205 66.120 ;
        RECT 40.735 66.090 41.385 66.120 ;
        RECT 36.770 65.835 37.000 65.980 ;
        RECT 38.410 65.835 38.640 65.980 ;
        RECT 40.345 65.835 40.575 65.980 ;
        RECT 41.545 65.835 41.775 65.980 ;
        RECT 41.980 65.835 42.270 66.710 ;
        RECT 36.770 65.665 42.270 65.835 ;
        RECT 36.315 65.380 36.615 65.635 ;
        RECT 36.770 65.520 37.000 65.665 ;
        RECT 38.410 65.520 38.640 65.665 ;
        RECT 40.345 65.520 40.575 65.665 ;
        RECT 41.545 65.520 41.775 65.665 ;
        RECT 37.205 65.380 38.205 65.410 ;
        RECT 40.735 65.380 41.385 65.410 ;
        RECT 41.980 65.380 42.270 65.665 ;
        RECT 43.030 66.710 44.935 66.880 ;
        RECT 47.425 66.775 48.985 66.880 ;
        RECT 49.740 66.880 50.030 68.210 ;
        RECT 50.625 68.180 51.625 68.210 ;
        RECT 51.870 67.950 52.130 68.270 ;
        RECT 54.135 68.210 55.690 68.380 ;
        RECT 56.445 68.380 56.745 68.635 ;
        RECT 56.900 68.520 57.130 68.665 ;
        RECT 58.540 68.520 58.770 68.665 ;
        RECT 59.470 68.590 59.730 68.665 ;
        RECT 60.475 68.520 60.705 68.665 ;
        RECT 61.675 68.520 61.905 68.665 ;
        RECT 57.335 68.380 58.335 68.410 ;
        RECT 60.865 68.380 61.515 68.410 ;
        RECT 62.110 68.380 62.400 69.710 ;
        RECT 63.160 69.710 65.065 69.880 ;
        RECT 67.555 69.775 69.115 69.880 ;
        RECT 69.870 69.880 70.160 71.275 ;
        RECT 70.735 71.210 71.775 71.380 ;
        RECT 74.265 71.210 75.820 71.380 ;
        RECT 76.575 71.275 76.875 71.635 ;
        RECT 77.030 71.520 77.260 71.665 ;
        RECT 77.865 71.590 78.125 71.665 ;
        RECT 78.670 71.520 78.900 71.665 ;
        RECT 80.605 71.520 80.835 71.665 ;
        RECT 81.805 71.520 82.035 71.665 ;
        RECT 77.465 71.380 78.465 71.410 ;
        RECT 80.995 71.380 81.645 71.410 ;
        RECT 82.240 71.380 82.530 72.710 ;
        RECT 83.290 71.635 83.580 74.210 ;
        RECT 84.175 74.180 85.175 74.210 ;
        RECT 87.705 74.180 88.355 74.210 ;
        RECT 84.175 73.790 85.175 73.820 ;
        RECT 86.310 73.790 86.570 73.865 ;
        RECT 87.705 73.790 88.355 73.820 ;
        RECT 84.155 73.620 88.375 73.790 ;
        RECT 84.175 73.590 85.175 73.620 ;
        RECT 86.310 73.545 86.570 73.620 ;
        RECT 87.705 73.590 88.355 73.620 ;
        RECT 83.740 73.335 83.970 73.480 ;
        RECT 84.155 73.335 84.415 73.410 ;
        RECT 85.380 73.335 85.610 73.480 ;
        RECT 87.315 73.335 87.545 73.480 ;
        RECT 88.515 73.335 88.745 73.480 ;
        RECT 83.740 73.165 88.745 73.335 ;
        RECT 83.740 73.020 83.970 73.165 ;
        RECT 84.155 73.090 84.415 73.165 ;
        RECT 85.380 73.020 85.610 73.165 ;
        RECT 87.315 73.020 87.545 73.165 ;
        RECT 88.515 73.020 88.745 73.165 ;
        RECT 88.950 73.135 89.240 74.210 ;
        RECT 90.000 74.210 91.905 74.275 ;
        RECT 94.395 74.210 95.950 74.380 ;
        RECT 96.705 74.380 97.005 74.635 ;
        RECT 97.160 74.520 97.390 74.665 ;
        RECT 98.800 74.590 99.095 74.665 ;
        RECT 98.800 74.520 99.030 74.590 ;
        RECT 100.735 74.520 100.965 74.665 ;
        RECT 101.935 74.520 102.165 74.665 ;
        RECT 97.595 74.380 98.595 74.410 ;
        RECT 101.125 74.380 101.775 74.410 ;
        RECT 102.370 74.380 102.660 75.710 ;
        RECT 96.705 74.275 98.615 74.380 ;
        RECT 84.175 72.880 85.175 72.910 ;
        RECT 87.705 72.880 88.355 72.910 ;
        RECT 88.945 72.880 89.245 73.135 ;
        RECT 84.155 72.710 85.195 72.880 ;
        RECT 87.685 72.775 89.245 72.880 ;
        RECT 87.685 72.710 89.240 72.775 ;
        RECT 84.175 72.680 85.175 72.710 ;
        RECT 87.705 72.680 88.355 72.710 ;
        RECT 84.590 72.320 84.760 72.680 ;
        RECT 84.175 72.290 85.175 72.320 ;
        RECT 86.310 72.290 86.570 72.365 ;
        RECT 87.705 72.290 88.355 72.320 ;
        RECT 84.155 72.120 85.195 72.290 ;
        RECT 86.310 72.120 88.375 72.290 ;
        RECT 84.175 72.090 85.175 72.120 ;
        RECT 86.310 72.045 86.570 72.120 ;
        RECT 87.705 72.090 88.355 72.120 ;
        RECT 83.740 71.835 83.970 71.980 ;
        RECT 84.575 71.835 84.835 71.910 ;
        RECT 85.380 71.835 85.610 71.980 ;
        RECT 87.315 71.835 87.545 71.980 ;
        RECT 88.515 71.835 88.745 71.980 ;
        RECT 83.740 71.665 88.745 71.835 ;
        RECT 70.755 71.180 71.755 71.210 ;
        RECT 74.285 71.180 74.935 71.210 ;
        RECT 71.170 70.820 71.340 71.180 ;
        RECT 70.755 70.790 71.755 70.820 ;
        RECT 72.890 70.790 73.150 70.865 ;
        RECT 74.285 70.790 74.935 70.820 ;
        RECT 70.735 70.620 71.775 70.790 ;
        RECT 72.890 70.620 74.955 70.790 ;
        RECT 70.755 70.590 71.755 70.620 ;
        RECT 72.890 70.545 73.150 70.620 ;
        RECT 74.285 70.590 74.935 70.620 ;
        RECT 70.320 70.335 70.550 70.480 ;
        RECT 71.960 70.410 72.190 70.480 ;
        RECT 71.960 70.335 72.255 70.410 ;
        RECT 73.895 70.335 74.125 70.480 ;
        RECT 75.095 70.335 75.325 70.480 ;
        RECT 70.320 70.165 75.325 70.335 ;
        RECT 70.320 70.020 70.550 70.165 ;
        RECT 71.960 70.090 72.255 70.165 ;
        RECT 71.960 70.020 72.190 70.090 ;
        RECT 73.895 70.020 74.125 70.165 ;
        RECT 75.095 70.020 75.325 70.165 ;
        RECT 75.530 70.135 75.820 71.210 ;
        RECT 70.755 69.880 71.755 69.910 ;
        RECT 74.285 69.880 74.935 69.910 ;
        RECT 75.525 69.880 75.825 70.135 ;
        RECT 67.555 69.710 69.110 69.775 ;
        RECT 63.160 68.635 63.450 69.710 ;
        RECT 64.045 69.680 65.045 69.710 ;
        RECT 67.575 69.680 68.225 69.710 ;
        RECT 67.985 69.320 68.245 69.365 ;
        RECT 64.045 69.290 65.045 69.320 ;
        RECT 67.575 69.290 68.245 69.320 ;
        RECT 64.025 69.120 68.245 69.290 ;
        RECT 64.045 69.090 65.045 69.120 ;
        RECT 67.575 69.090 68.245 69.120 ;
        RECT 67.985 69.045 68.245 69.090 ;
        RECT 63.610 68.835 63.840 68.980 ;
        RECT 65.250 68.835 65.480 68.980 ;
        RECT 66.180 68.835 66.440 68.910 ;
        RECT 67.185 68.835 67.415 68.980 ;
        RECT 68.385 68.835 68.615 68.980 ;
        RECT 63.610 68.665 68.615 68.835 ;
        RECT 56.445 68.275 58.355 68.380 ;
        RECT 54.155 68.180 54.805 68.210 ;
        RECT 50.625 67.790 51.625 67.820 ;
        RECT 51.915 67.790 52.085 67.950 ;
        RECT 52.760 67.790 53.020 67.865 ;
        RECT 54.155 67.790 54.805 67.820 ;
        RECT 50.605 67.620 54.825 67.790 ;
        RECT 50.625 67.590 51.625 67.620 ;
        RECT 52.760 67.545 53.020 67.620 ;
        RECT 54.155 67.590 54.805 67.620 ;
        RECT 50.190 67.335 50.420 67.480 ;
        RECT 51.830 67.335 52.060 67.480 ;
        RECT 52.730 67.335 53.050 67.380 ;
        RECT 53.765 67.335 53.995 67.480 ;
        RECT 54.965 67.335 55.195 67.480 ;
        RECT 50.190 67.165 55.195 67.335 ;
        RECT 50.190 67.020 50.420 67.165 ;
        RECT 51.830 67.020 52.060 67.165 ;
        RECT 52.730 67.120 53.050 67.165 ;
        RECT 53.765 67.020 53.995 67.165 ;
        RECT 54.965 67.020 55.195 67.165 ;
        RECT 55.400 67.135 55.690 68.210 ;
        RECT 56.450 68.210 58.355 68.275 ;
        RECT 60.845 68.210 62.400 68.380 ;
        RECT 63.155 68.380 63.455 68.635 ;
        RECT 63.610 68.520 63.840 68.665 ;
        RECT 65.250 68.520 65.480 68.665 ;
        RECT 66.180 68.590 66.440 68.665 ;
        RECT 67.185 68.520 67.415 68.665 ;
        RECT 68.385 68.520 68.615 68.665 ;
        RECT 64.045 68.380 65.045 68.410 ;
        RECT 67.575 68.380 68.225 68.410 ;
        RECT 68.820 68.380 69.110 69.710 ;
        RECT 69.870 69.710 71.775 69.880 ;
        RECT 74.265 69.775 75.825 69.880 ;
        RECT 76.580 69.880 76.870 71.275 ;
        RECT 77.445 71.210 78.485 71.380 ;
        RECT 80.975 71.210 82.530 71.380 ;
        RECT 83.285 71.275 83.585 71.635 ;
        RECT 83.740 71.520 83.970 71.665 ;
        RECT 84.575 71.590 84.835 71.665 ;
        RECT 85.380 71.520 85.610 71.665 ;
        RECT 87.315 71.520 87.545 71.665 ;
        RECT 88.515 71.520 88.745 71.665 ;
        RECT 84.175 71.380 85.175 71.410 ;
        RECT 87.705 71.380 88.355 71.410 ;
        RECT 88.950 71.380 89.240 72.710 ;
        RECT 90.000 71.635 90.290 74.210 ;
        RECT 90.885 74.180 91.885 74.210 ;
        RECT 94.415 74.180 95.065 74.210 ;
        RECT 90.885 73.790 91.885 73.820 ;
        RECT 93.020 73.790 93.280 73.865 ;
        RECT 94.415 73.790 95.065 73.820 ;
        RECT 90.865 73.620 95.085 73.790 ;
        RECT 90.885 73.590 91.885 73.620 ;
        RECT 93.020 73.545 93.280 73.620 ;
        RECT 94.415 73.590 95.065 73.620 ;
        RECT 90.450 73.335 90.680 73.480 ;
        RECT 90.865 73.335 91.125 73.410 ;
        RECT 92.090 73.335 92.320 73.480 ;
        RECT 94.025 73.335 94.255 73.480 ;
        RECT 95.225 73.335 95.455 73.480 ;
        RECT 90.450 73.165 95.455 73.335 ;
        RECT 90.450 73.020 90.680 73.165 ;
        RECT 90.865 73.090 91.125 73.165 ;
        RECT 92.090 73.020 92.320 73.165 ;
        RECT 94.025 73.020 94.255 73.165 ;
        RECT 95.225 73.020 95.455 73.165 ;
        RECT 95.660 73.135 95.950 74.210 ;
        RECT 96.710 74.210 98.615 74.275 ;
        RECT 101.105 74.210 102.660 74.380 ;
        RECT 90.885 72.880 91.885 72.910 ;
        RECT 94.415 72.880 95.065 72.910 ;
        RECT 95.655 72.880 95.955 73.135 ;
        RECT 90.865 72.710 91.905 72.880 ;
        RECT 94.395 72.775 95.955 72.880 ;
        RECT 94.395 72.710 95.950 72.775 ;
        RECT 90.885 72.680 91.885 72.710 ;
        RECT 94.415 72.680 95.065 72.710 ;
        RECT 91.300 72.320 91.470 72.680 ;
        RECT 90.885 72.290 91.885 72.320 ;
        RECT 93.020 72.290 93.280 72.365 ;
        RECT 94.415 72.290 95.065 72.320 ;
        RECT 90.865 72.120 91.905 72.290 ;
        RECT 93.020 72.120 95.085 72.290 ;
        RECT 90.885 72.090 91.885 72.120 ;
        RECT 93.020 72.045 93.280 72.120 ;
        RECT 94.415 72.090 95.065 72.120 ;
        RECT 90.450 71.835 90.680 71.980 ;
        RECT 91.285 71.835 91.545 71.910 ;
        RECT 92.090 71.835 92.320 71.980 ;
        RECT 94.025 71.835 94.255 71.980 ;
        RECT 95.225 71.835 95.455 71.980 ;
        RECT 90.450 71.665 95.455 71.835 ;
        RECT 77.465 71.180 78.465 71.210 ;
        RECT 80.995 71.180 81.645 71.210 ;
        RECT 77.880 70.820 78.050 71.180 ;
        RECT 77.465 70.790 78.465 70.820 ;
        RECT 79.600 70.790 79.860 70.865 ;
        RECT 80.995 70.790 81.645 70.820 ;
        RECT 77.445 70.620 78.485 70.790 ;
        RECT 79.600 70.620 81.665 70.790 ;
        RECT 77.465 70.590 78.465 70.620 ;
        RECT 79.600 70.545 79.860 70.620 ;
        RECT 80.995 70.590 81.645 70.620 ;
        RECT 77.030 70.335 77.260 70.480 ;
        RECT 78.670 70.410 78.900 70.480 ;
        RECT 78.670 70.335 78.965 70.410 ;
        RECT 80.605 70.335 80.835 70.480 ;
        RECT 81.805 70.335 82.035 70.480 ;
        RECT 77.030 70.165 82.035 70.335 ;
        RECT 77.030 70.020 77.260 70.165 ;
        RECT 78.670 70.090 78.965 70.165 ;
        RECT 78.670 70.020 78.900 70.090 ;
        RECT 80.605 70.020 80.835 70.165 ;
        RECT 81.805 70.020 82.035 70.165 ;
        RECT 82.240 70.135 82.530 71.210 ;
        RECT 77.465 69.880 78.465 69.910 ;
        RECT 80.995 69.880 81.645 69.910 ;
        RECT 82.235 69.880 82.535 70.135 ;
        RECT 74.265 69.710 75.820 69.775 ;
        RECT 69.870 68.635 70.160 69.710 ;
        RECT 70.755 69.680 71.755 69.710 ;
        RECT 74.285 69.680 74.935 69.710 ;
        RECT 71.155 69.320 71.415 69.365 ;
        RECT 70.755 69.290 71.755 69.320 ;
        RECT 74.285 69.290 74.935 69.320 ;
        RECT 70.735 69.120 74.955 69.290 ;
        RECT 70.755 69.090 71.755 69.120 ;
        RECT 74.285 69.090 74.935 69.120 ;
        RECT 71.155 69.045 71.415 69.090 ;
        RECT 70.320 68.835 70.550 68.980 ;
        RECT 71.960 68.835 72.190 68.980 ;
        RECT 72.890 68.835 73.150 68.910 ;
        RECT 73.895 68.835 74.125 68.980 ;
        RECT 75.095 68.835 75.325 68.980 ;
        RECT 70.320 68.665 75.325 68.835 ;
        RECT 63.155 68.275 65.065 68.380 ;
        RECT 50.625 66.880 51.625 66.910 ;
        RECT 54.155 66.880 54.805 66.910 ;
        RECT 55.395 66.880 55.695 67.135 ;
        RECT 47.425 66.710 48.980 66.775 ;
        RECT 43.030 65.635 43.320 66.710 ;
        RECT 43.915 66.680 44.915 66.710 ;
        RECT 47.445 66.680 48.095 66.710 ;
        RECT 43.895 66.320 44.155 66.365 ;
        RECT 43.895 66.290 44.915 66.320 ;
        RECT 47.445 66.290 48.095 66.320 ;
        RECT 43.895 66.120 48.115 66.290 ;
        RECT 43.895 66.090 44.915 66.120 ;
        RECT 47.445 66.090 48.095 66.120 ;
        RECT 43.895 66.045 44.155 66.090 ;
        RECT 43.480 65.835 43.710 65.980 ;
        RECT 45.120 65.835 45.350 65.980 ;
        RECT 47.055 65.835 47.285 65.980 ;
        RECT 47.855 65.835 48.115 65.910 ;
        RECT 48.255 65.835 48.485 65.980 ;
        RECT 43.480 65.665 48.485 65.835 ;
        RECT 36.315 65.275 38.225 65.380 ;
        RECT 36.320 65.210 38.225 65.275 ;
        RECT 40.715 65.210 42.270 65.380 ;
        RECT 43.025 65.380 43.325 65.635 ;
        RECT 43.480 65.520 43.710 65.665 ;
        RECT 45.120 65.520 45.350 65.665 ;
        RECT 47.055 65.520 47.285 65.665 ;
        RECT 47.855 65.590 48.115 65.665 ;
        RECT 48.255 65.520 48.485 65.665 ;
        RECT 43.915 65.380 44.915 65.410 ;
        RECT 47.445 65.380 48.095 65.410 ;
        RECT 48.690 65.380 48.980 66.710 ;
        RECT 49.740 66.710 51.645 66.880 ;
        RECT 54.135 66.775 55.695 66.880 ;
        RECT 56.450 66.880 56.740 68.210 ;
        RECT 57.335 68.180 58.335 68.210 ;
        RECT 60.865 68.180 61.515 68.210 ;
        RECT 58.155 67.820 58.415 67.865 ;
        RECT 57.335 67.790 58.415 67.820 ;
        RECT 59.470 67.790 59.730 67.865 ;
        RECT 60.865 67.790 61.515 67.820 ;
        RECT 57.315 67.620 61.535 67.790 ;
        RECT 57.335 67.590 58.415 67.620 ;
        RECT 58.155 67.545 58.415 67.590 ;
        RECT 59.470 67.545 59.730 67.620 ;
        RECT 60.865 67.590 61.515 67.620 ;
        RECT 56.900 67.335 57.130 67.480 ;
        RECT 58.540 67.335 58.770 67.480 ;
        RECT 59.440 67.335 59.760 67.380 ;
        RECT 60.475 67.335 60.705 67.480 ;
        RECT 61.675 67.335 61.905 67.480 ;
        RECT 56.900 67.165 61.905 67.335 ;
        RECT 56.900 67.020 57.130 67.165 ;
        RECT 58.540 67.020 58.770 67.165 ;
        RECT 59.440 67.120 59.760 67.165 ;
        RECT 60.475 67.020 60.705 67.165 ;
        RECT 61.675 67.020 61.905 67.165 ;
        RECT 62.110 67.135 62.400 68.210 ;
        RECT 63.160 68.210 65.065 68.275 ;
        RECT 57.335 66.880 58.335 66.910 ;
        RECT 60.865 66.880 61.515 66.910 ;
        RECT 62.105 66.880 62.405 67.135 ;
        RECT 54.135 66.710 55.690 66.775 ;
        RECT 49.740 65.635 50.030 66.710 ;
        RECT 50.625 66.680 51.625 66.710 ;
        RECT 54.155 66.680 54.805 66.710 ;
        RECT 50.625 66.290 51.625 66.320 ;
        RECT 54.155 66.290 54.805 66.320 ;
        RECT 50.605 66.120 54.825 66.290 ;
        RECT 50.625 66.090 51.625 66.120 ;
        RECT 54.155 66.090 54.805 66.120 ;
        RECT 50.190 65.835 50.420 65.980 ;
        RECT 51.830 65.835 52.060 65.980 ;
        RECT 53.765 65.835 53.995 65.980 ;
        RECT 54.965 65.835 55.195 65.980 ;
        RECT 55.400 65.835 55.690 66.710 ;
        RECT 50.190 65.665 55.690 65.835 ;
        RECT 43.025 65.275 44.935 65.380 ;
        RECT 36.320 65.000 36.610 65.210 ;
        RECT 37.205 65.180 38.205 65.210 ;
        RECT 40.735 65.180 41.385 65.210 ;
        RECT 41.980 65.000 42.270 65.210 ;
        RECT 43.030 65.210 44.935 65.275 ;
        RECT 47.425 65.210 48.980 65.380 ;
        RECT 49.735 65.380 50.035 65.635 ;
        RECT 50.190 65.520 50.420 65.665 ;
        RECT 51.830 65.520 52.060 65.665 ;
        RECT 53.765 65.520 53.995 65.665 ;
        RECT 54.965 65.520 55.195 65.665 ;
        RECT 50.625 65.380 51.625 65.410 ;
        RECT 54.155 65.380 54.805 65.410 ;
        RECT 55.400 65.380 55.690 65.665 ;
        RECT 56.450 66.710 58.355 66.880 ;
        RECT 60.845 66.775 62.405 66.880 ;
        RECT 63.160 66.880 63.450 68.210 ;
        RECT 64.045 68.180 65.045 68.210 ;
        RECT 65.290 67.950 65.550 68.270 ;
        RECT 67.555 68.210 69.110 68.380 ;
        RECT 69.865 68.380 70.165 68.635 ;
        RECT 70.320 68.520 70.550 68.665 ;
        RECT 71.960 68.520 72.190 68.665 ;
        RECT 72.890 68.590 73.150 68.665 ;
        RECT 73.895 68.520 74.125 68.665 ;
        RECT 75.095 68.520 75.325 68.665 ;
        RECT 70.755 68.380 71.755 68.410 ;
        RECT 74.285 68.380 74.935 68.410 ;
        RECT 75.530 68.380 75.820 69.710 ;
        RECT 76.580 69.710 78.485 69.880 ;
        RECT 80.975 69.775 82.535 69.880 ;
        RECT 83.290 69.880 83.580 71.275 ;
        RECT 84.155 71.210 85.195 71.380 ;
        RECT 87.685 71.210 89.240 71.380 ;
        RECT 89.995 71.275 90.295 71.635 ;
        RECT 90.450 71.520 90.680 71.665 ;
        RECT 91.285 71.590 91.545 71.665 ;
        RECT 92.090 71.520 92.320 71.665 ;
        RECT 94.025 71.520 94.255 71.665 ;
        RECT 95.225 71.520 95.455 71.665 ;
        RECT 90.885 71.380 91.885 71.410 ;
        RECT 94.415 71.380 95.065 71.410 ;
        RECT 95.660 71.380 95.950 72.710 ;
        RECT 96.710 71.635 97.000 74.210 ;
        RECT 97.595 74.180 98.595 74.210 ;
        RECT 101.125 74.180 101.775 74.210 ;
        RECT 97.595 73.790 98.595 73.820 ;
        RECT 99.730 73.790 99.990 73.865 ;
        RECT 101.125 73.790 101.775 73.820 ;
        RECT 97.575 73.620 101.795 73.790 ;
        RECT 97.595 73.590 98.595 73.620 ;
        RECT 99.730 73.545 99.990 73.620 ;
        RECT 101.125 73.590 101.775 73.620 ;
        RECT 97.160 73.335 97.390 73.480 ;
        RECT 97.575 73.335 97.835 73.410 ;
        RECT 98.800 73.335 99.030 73.480 ;
        RECT 100.735 73.335 100.965 73.480 ;
        RECT 101.935 73.335 102.165 73.480 ;
        RECT 97.160 73.165 102.165 73.335 ;
        RECT 97.160 73.020 97.390 73.165 ;
        RECT 97.575 73.090 97.835 73.165 ;
        RECT 98.800 73.020 99.030 73.165 ;
        RECT 100.735 73.020 100.965 73.165 ;
        RECT 101.935 73.020 102.165 73.165 ;
        RECT 102.370 73.135 102.660 74.210 ;
        RECT 97.595 72.880 98.595 72.910 ;
        RECT 101.125 72.880 101.775 72.910 ;
        RECT 102.365 72.880 102.665 73.135 ;
        RECT 97.575 72.710 98.615 72.880 ;
        RECT 101.105 72.775 102.665 72.880 ;
        RECT 101.105 72.710 102.660 72.775 ;
        RECT 97.595 72.680 98.595 72.710 ;
        RECT 101.125 72.680 101.775 72.710 ;
        RECT 98.010 72.320 98.180 72.680 ;
        RECT 97.595 72.290 98.595 72.320 ;
        RECT 99.730 72.290 99.990 72.365 ;
        RECT 101.125 72.290 101.775 72.320 ;
        RECT 97.575 72.120 98.615 72.290 ;
        RECT 99.730 72.120 101.795 72.290 ;
        RECT 97.595 72.090 98.595 72.120 ;
        RECT 99.730 72.045 99.990 72.120 ;
        RECT 101.125 72.090 101.775 72.120 ;
        RECT 97.160 71.835 97.390 71.980 ;
        RECT 97.995 71.835 98.255 71.910 ;
        RECT 98.800 71.835 99.030 71.980 ;
        RECT 100.735 71.835 100.965 71.980 ;
        RECT 101.935 71.835 102.165 71.980 ;
        RECT 97.160 71.665 102.165 71.835 ;
        RECT 84.175 71.180 85.175 71.210 ;
        RECT 87.705 71.180 88.355 71.210 ;
        RECT 84.590 70.820 84.760 71.180 ;
        RECT 84.175 70.790 85.175 70.820 ;
        RECT 86.310 70.790 86.570 70.865 ;
        RECT 87.705 70.790 88.355 70.820 ;
        RECT 84.155 70.620 85.195 70.790 ;
        RECT 86.310 70.620 88.375 70.790 ;
        RECT 84.175 70.590 85.175 70.620 ;
        RECT 86.310 70.545 86.570 70.620 ;
        RECT 87.705 70.590 88.355 70.620 ;
        RECT 83.740 70.335 83.970 70.480 ;
        RECT 85.380 70.410 85.610 70.480 ;
        RECT 85.380 70.335 85.675 70.410 ;
        RECT 87.315 70.335 87.545 70.480 ;
        RECT 88.515 70.335 88.745 70.480 ;
        RECT 83.740 70.165 88.745 70.335 ;
        RECT 83.740 70.020 83.970 70.165 ;
        RECT 85.380 70.090 85.675 70.165 ;
        RECT 85.380 70.020 85.610 70.090 ;
        RECT 87.315 70.020 87.545 70.165 ;
        RECT 88.515 70.020 88.745 70.165 ;
        RECT 88.950 70.135 89.240 71.210 ;
        RECT 84.175 69.880 85.175 69.910 ;
        RECT 87.705 69.880 88.355 69.910 ;
        RECT 88.945 69.880 89.245 70.135 ;
        RECT 80.975 69.710 82.530 69.775 ;
        RECT 76.580 68.635 76.870 69.710 ;
        RECT 77.465 69.680 78.465 69.710 ;
        RECT 80.995 69.680 81.645 69.710 ;
        RECT 81.405 69.320 81.665 69.365 ;
        RECT 77.465 69.290 78.465 69.320 ;
        RECT 80.995 69.290 81.665 69.320 ;
        RECT 77.445 69.120 81.665 69.290 ;
        RECT 77.465 69.090 78.465 69.120 ;
        RECT 80.995 69.090 81.665 69.120 ;
        RECT 81.405 69.045 81.665 69.090 ;
        RECT 77.030 68.835 77.260 68.980 ;
        RECT 78.670 68.835 78.900 68.980 ;
        RECT 79.600 68.835 79.860 68.910 ;
        RECT 80.605 68.835 80.835 68.980 ;
        RECT 81.805 68.835 82.035 68.980 ;
        RECT 77.030 68.665 82.035 68.835 ;
        RECT 69.865 68.275 71.775 68.380 ;
        RECT 67.575 68.180 68.225 68.210 ;
        RECT 64.045 67.790 65.045 67.820 ;
        RECT 65.335 67.790 65.505 67.950 ;
        RECT 66.180 67.790 66.440 67.865 ;
        RECT 67.575 67.790 68.225 67.820 ;
        RECT 64.025 67.620 68.245 67.790 ;
        RECT 64.045 67.590 65.045 67.620 ;
        RECT 66.180 67.545 66.440 67.620 ;
        RECT 67.575 67.590 68.225 67.620 ;
        RECT 63.610 67.335 63.840 67.480 ;
        RECT 65.250 67.335 65.480 67.480 ;
        RECT 66.150 67.335 66.470 67.380 ;
        RECT 67.185 67.335 67.415 67.480 ;
        RECT 68.385 67.335 68.615 67.480 ;
        RECT 63.610 67.165 68.615 67.335 ;
        RECT 63.610 67.020 63.840 67.165 ;
        RECT 65.250 67.020 65.480 67.165 ;
        RECT 66.150 67.120 66.470 67.165 ;
        RECT 67.185 67.020 67.415 67.165 ;
        RECT 68.385 67.020 68.615 67.165 ;
        RECT 68.820 67.135 69.110 68.210 ;
        RECT 69.870 68.210 71.775 68.275 ;
        RECT 74.265 68.210 75.820 68.380 ;
        RECT 76.575 68.380 76.875 68.635 ;
        RECT 77.030 68.520 77.260 68.665 ;
        RECT 78.670 68.520 78.900 68.665 ;
        RECT 79.600 68.590 79.860 68.665 ;
        RECT 80.605 68.520 80.835 68.665 ;
        RECT 81.805 68.520 82.035 68.665 ;
        RECT 77.465 68.380 78.465 68.410 ;
        RECT 80.995 68.380 81.645 68.410 ;
        RECT 82.240 68.380 82.530 69.710 ;
        RECT 83.290 69.710 85.195 69.880 ;
        RECT 87.685 69.775 89.245 69.880 ;
        RECT 90.000 69.880 90.290 71.275 ;
        RECT 90.865 71.210 91.905 71.380 ;
        RECT 94.395 71.210 95.950 71.380 ;
        RECT 96.705 71.275 97.005 71.635 ;
        RECT 97.160 71.520 97.390 71.665 ;
        RECT 97.995 71.590 98.255 71.665 ;
        RECT 98.800 71.520 99.030 71.665 ;
        RECT 100.735 71.520 100.965 71.665 ;
        RECT 101.935 71.520 102.165 71.665 ;
        RECT 97.595 71.380 98.595 71.410 ;
        RECT 101.125 71.380 101.775 71.410 ;
        RECT 102.370 71.380 102.660 72.710 ;
        RECT 90.885 71.180 91.885 71.210 ;
        RECT 94.415 71.180 95.065 71.210 ;
        RECT 91.300 70.820 91.470 71.180 ;
        RECT 90.885 70.790 91.885 70.820 ;
        RECT 93.020 70.790 93.280 70.865 ;
        RECT 94.415 70.790 95.065 70.820 ;
        RECT 90.865 70.620 91.905 70.790 ;
        RECT 93.020 70.620 95.085 70.790 ;
        RECT 90.885 70.590 91.885 70.620 ;
        RECT 93.020 70.545 93.280 70.620 ;
        RECT 94.415 70.590 95.065 70.620 ;
        RECT 90.450 70.335 90.680 70.480 ;
        RECT 92.090 70.410 92.320 70.480 ;
        RECT 92.090 70.335 92.385 70.410 ;
        RECT 94.025 70.335 94.255 70.480 ;
        RECT 95.225 70.335 95.455 70.480 ;
        RECT 90.450 70.165 95.455 70.335 ;
        RECT 90.450 70.020 90.680 70.165 ;
        RECT 92.090 70.090 92.385 70.165 ;
        RECT 92.090 70.020 92.320 70.090 ;
        RECT 94.025 70.020 94.255 70.165 ;
        RECT 95.225 70.020 95.455 70.165 ;
        RECT 95.660 70.135 95.950 71.210 ;
        RECT 90.885 69.880 91.885 69.910 ;
        RECT 94.415 69.880 95.065 69.910 ;
        RECT 95.655 69.880 95.955 70.135 ;
        RECT 87.685 69.710 89.240 69.775 ;
        RECT 83.290 68.635 83.580 69.710 ;
        RECT 84.175 69.680 85.175 69.710 ;
        RECT 87.705 69.680 88.355 69.710 ;
        RECT 84.575 69.320 84.835 69.365 ;
        RECT 84.175 69.290 85.175 69.320 ;
        RECT 87.705 69.290 88.355 69.320 ;
        RECT 84.155 69.120 88.375 69.290 ;
        RECT 84.175 69.090 85.175 69.120 ;
        RECT 87.705 69.090 88.355 69.120 ;
        RECT 84.575 69.045 84.835 69.090 ;
        RECT 83.740 68.835 83.970 68.980 ;
        RECT 85.380 68.835 85.610 68.980 ;
        RECT 86.310 68.835 86.570 68.910 ;
        RECT 87.315 68.835 87.545 68.980 ;
        RECT 88.515 68.835 88.745 68.980 ;
        RECT 83.740 68.665 88.745 68.835 ;
        RECT 76.575 68.275 78.485 68.380 ;
        RECT 64.045 66.880 65.045 66.910 ;
        RECT 67.575 66.880 68.225 66.910 ;
        RECT 68.815 66.880 69.115 67.135 ;
        RECT 60.845 66.710 62.400 66.775 ;
        RECT 56.450 65.635 56.740 66.710 ;
        RECT 57.335 66.680 58.335 66.710 ;
        RECT 60.865 66.680 61.515 66.710 ;
        RECT 57.315 66.320 57.575 66.365 ;
        RECT 57.315 66.290 58.335 66.320 ;
        RECT 60.865 66.290 61.515 66.320 ;
        RECT 57.315 66.120 61.535 66.290 ;
        RECT 57.315 66.090 58.335 66.120 ;
        RECT 60.865 66.090 61.515 66.120 ;
        RECT 57.315 66.045 57.575 66.090 ;
        RECT 56.900 65.835 57.130 65.980 ;
        RECT 58.540 65.835 58.770 65.980 ;
        RECT 60.475 65.835 60.705 65.980 ;
        RECT 61.275 65.835 61.535 65.910 ;
        RECT 61.675 65.835 61.905 65.980 ;
        RECT 56.900 65.665 61.905 65.835 ;
        RECT 49.735 65.275 51.645 65.380 ;
        RECT 43.030 65.000 43.320 65.210 ;
        RECT 43.915 65.180 44.915 65.210 ;
        RECT 47.445 65.180 48.095 65.210 ;
        RECT 48.690 65.000 48.980 65.210 ;
        RECT 49.740 65.210 51.645 65.275 ;
        RECT 54.135 65.210 55.690 65.380 ;
        RECT 56.445 65.380 56.745 65.635 ;
        RECT 56.900 65.520 57.130 65.665 ;
        RECT 58.540 65.520 58.770 65.665 ;
        RECT 60.475 65.520 60.705 65.665 ;
        RECT 61.275 65.590 61.535 65.665 ;
        RECT 61.675 65.520 61.905 65.665 ;
        RECT 57.335 65.380 58.335 65.410 ;
        RECT 60.865 65.380 61.515 65.410 ;
        RECT 62.110 65.380 62.400 66.710 ;
        RECT 63.160 66.710 65.065 66.880 ;
        RECT 67.555 66.775 69.115 66.880 ;
        RECT 69.870 66.880 70.160 68.210 ;
        RECT 70.755 68.180 71.755 68.210 ;
        RECT 74.285 68.180 74.935 68.210 ;
        RECT 71.575 67.820 71.835 67.865 ;
        RECT 70.755 67.790 71.835 67.820 ;
        RECT 72.890 67.790 73.150 67.865 ;
        RECT 74.285 67.790 74.935 67.820 ;
        RECT 70.735 67.620 74.955 67.790 ;
        RECT 70.755 67.590 71.835 67.620 ;
        RECT 71.575 67.545 71.835 67.590 ;
        RECT 72.890 67.545 73.150 67.620 ;
        RECT 74.285 67.590 74.935 67.620 ;
        RECT 70.320 67.335 70.550 67.480 ;
        RECT 71.960 67.335 72.190 67.480 ;
        RECT 72.860 67.335 73.180 67.380 ;
        RECT 73.895 67.335 74.125 67.480 ;
        RECT 75.095 67.335 75.325 67.480 ;
        RECT 70.320 67.165 75.325 67.335 ;
        RECT 70.320 67.020 70.550 67.165 ;
        RECT 71.960 67.020 72.190 67.165 ;
        RECT 72.860 67.120 73.180 67.165 ;
        RECT 73.895 67.020 74.125 67.165 ;
        RECT 75.095 67.020 75.325 67.165 ;
        RECT 75.530 67.135 75.820 68.210 ;
        RECT 76.580 68.210 78.485 68.275 ;
        RECT 70.755 66.880 71.755 66.910 ;
        RECT 74.285 66.880 74.935 66.910 ;
        RECT 75.525 66.880 75.825 67.135 ;
        RECT 67.555 66.710 69.110 66.775 ;
        RECT 63.160 65.635 63.450 66.710 ;
        RECT 64.045 66.680 65.045 66.710 ;
        RECT 67.575 66.680 68.225 66.710 ;
        RECT 64.045 66.290 65.045 66.320 ;
        RECT 67.575 66.290 68.225 66.320 ;
        RECT 64.025 66.120 68.245 66.290 ;
        RECT 64.045 66.090 65.045 66.120 ;
        RECT 67.575 66.090 68.225 66.120 ;
        RECT 63.610 65.835 63.840 65.980 ;
        RECT 65.250 65.835 65.480 65.980 ;
        RECT 67.185 65.835 67.415 65.980 ;
        RECT 68.385 65.835 68.615 65.980 ;
        RECT 68.820 65.835 69.110 66.710 ;
        RECT 63.610 65.665 69.110 65.835 ;
        RECT 56.445 65.275 58.355 65.380 ;
        RECT 49.740 65.000 50.030 65.210 ;
        RECT 50.625 65.180 51.625 65.210 ;
        RECT 54.155 65.180 54.805 65.210 ;
        RECT 55.400 65.000 55.690 65.210 ;
        RECT 56.450 65.210 58.355 65.275 ;
        RECT 60.845 65.210 62.400 65.380 ;
        RECT 63.155 65.380 63.455 65.635 ;
        RECT 63.610 65.520 63.840 65.665 ;
        RECT 65.250 65.520 65.480 65.665 ;
        RECT 67.185 65.520 67.415 65.665 ;
        RECT 68.385 65.520 68.615 65.665 ;
        RECT 64.045 65.380 65.045 65.410 ;
        RECT 67.575 65.380 68.225 65.410 ;
        RECT 68.820 65.380 69.110 65.665 ;
        RECT 69.870 66.710 71.775 66.880 ;
        RECT 74.265 66.775 75.825 66.880 ;
        RECT 76.580 66.880 76.870 68.210 ;
        RECT 77.465 68.180 78.465 68.210 ;
        RECT 78.710 67.950 78.970 68.270 ;
        RECT 80.975 68.210 82.530 68.380 ;
        RECT 83.285 68.380 83.585 68.635 ;
        RECT 83.740 68.520 83.970 68.665 ;
        RECT 85.380 68.520 85.610 68.665 ;
        RECT 86.310 68.590 86.570 68.665 ;
        RECT 87.315 68.520 87.545 68.665 ;
        RECT 88.515 68.520 88.745 68.665 ;
        RECT 84.175 68.380 85.175 68.410 ;
        RECT 87.705 68.380 88.355 68.410 ;
        RECT 88.950 68.380 89.240 69.710 ;
        RECT 90.000 69.710 91.905 69.880 ;
        RECT 94.395 69.775 95.955 69.880 ;
        RECT 96.710 69.880 97.000 71.275 ;
        RECT 97.575 71.210 98.615 71.380 ;
        RECT 101.105 71.210 102.660 71.380 ;
        RECT 97.595 71.180 98.595 71.210 ;
        RECT 101.125 71.180 101.775 71.210 ;
        RECT 98.010 70.820 98.180 71.180 ;
        RECT 97.595 70.790 98.595 70.820 ;
        RECT 99.730 70.790 99.990 70.865 ;
        RECT 101.125 70.790 101.775 70.820 ;
        RECT 97.575 70.620 98.615 70.790 ;
        RECT 99.730 70.620 101.795 70.790 ;
        RECT 97.595 70.590 98.595 70.620 ;
        RECT 99.730 70.545 99.990 70.620 ;
        RECT 101.125 70.590 101.775 70.620 ;
        RECT 97.160 70.335 97.390 70.480 ;
        RECT 98.800 70.410 99.030 70.480 ;
        RECT 98.800 70.335 99.095 70.410 ;
        RECT 100.735 70.335 100.965 70.480 ;
        RECT 101.935 70.335 102.165 70.480 ;
        RECT 97.160 70.165 102.165 70.335 ;
        RECT 97.160 70.020 97.390 70.165 ;
        RECT 98.800 70.090 99.095 70.165 ;
        RECT 98.800 70.020 99.030 70.090 ;
        RECT 100.735 70.020 100.965 70.165 ;
        RECT 101.935 70.020 102.165 70.165 ;
        RECT 102.370 70.135 102.660 71.210 ;
        RECT 97.595 69.880 98.595 69.910 ;
        RECT 101.125 69.880 101.775 69.910 ;
        RECT 102.365 69.880 102.665 70.135 ;
        RECT 94.395 69.710 95.950 69.775 ;
        RECT 90.000 68.635 90.290 69.710 ;
        RECT 90.885 69.680 91.885 69.710 ;
        RECT 94.415 69.680 95.065 69.710 ;
        RECT 94.825 69.320 95.085 69.365 ;
        RECT 90.885 69.290 91.885 69.320 ;
        RECT 94.415 69.290 95.085 69.320 ;
        RECT 90.865 69.120 95.085 69.290 ;
        RECT 90.885 69.090 91.885 69.120 ;
        RECT 94.415 69.090 95.085 69.120 ;
        RECT 94.825 69.045 95.085 69.090 ;
        RECT 90.450 68.835 90.680 68.980 ;
        RECT 92.090 68.835 92.320 68.980 ;
        RECT 93.020 68.835 93.280 68.910 ;
        RECT 94.025 68.835 94.255 68.980 ;
        RECT 95.225 68.835 95.455 68.980 ;
        RECT 90.450 68.665 95.455 68.835 ;
        RECT 83.285 68.275 85.195 68.380 ;
        RECT 80.995 68.180 81.645 68.210 ;
        RECT 77.465 67.790 78.465 67.820 ;
        RECT 78.755 67.790 78.925 67.950 ;
        RECT 79.600 67.790 79.860 67.865 ;
        RECT 80.995 67.790 81.645 67.820 ;
        RECT 77.445 67.620 81.665 67.790 ;
        RECT 77.465 67.590 78.465 67.620 ;
        RECT 79.600 67.545 79.860 67.620 ;
        RECT 80.995 67.590 81.645 67.620 ;
        RECT 77.030 67.335 77.260 67.480 ;
        RECT 78.670 67.335 78.900 67.480 ;
        RECT 79.570 67.335 79.890 67.380 ;
        RECT 80.605 67.335 80.835 67.480 ;
        RECT 81.805 67.335 82.035 67.480 ;
        RECT 77.030 67.165 82.035 67.335 ;
        RECT 77.030 67.020 77.260 67.165 ;
        RECT 78.670 67.020 78.900 67.165 ;
        RECT 79.570 67.120 79.890 67.165 ;
        RECT 80.605 67.020 80.835 67.165 ;
        RECT 81.805 67.020 82.035 67.165 ;
        RECT 82.240 67.135 82.530 68.210 ;
        RECT 83.290 68.210 85.195 68.275 ;
        RECT 87.685 68.210 89.240 68.380 ;
        RECT 89.995 68.380 90.295 68.635 ;
        RECT 90.450 68.520 90.680 68.665 ;
        RECT 92.090 68.520 92.320 68.665 ;
        RECT 93.020 68.590 93.280 68.665 ;
        RECT 94.025 68.520 94.255 68.665 ;
        RECT 95.225 68.520 95.455 68.665 ;
        RECT 90.885 68.380 91.885 68.410 ;
        RECT 94.415 68.380 95.065 68.410 ;
        RECT 95.660 68.380 95.950 69.710 ;
        RECT 96.710 69.710 98.615 69.880 ;
        RECT 101.105 69.775 102.665 69.880 ;
        RECT 101.105 69.710 102.660 69.775 ;
        RECT 96.710 68.635 97.000 69.710 ;
        RECT 97.595 69.680 98.595 69.710 ;
        RECT 101.125 69.680 101.775 69.710 ;
        RECT 97.995 69.320 98.255 69.365 ;
        RECT 97.595 69.290 98.595 69.320 ;
        RECT 101.125 69.290 101.775 69.320 ;
        RECT 97.575 69.120 101.795 69.290 ;
        RECT 97.595 69.090 98.595 69.120 ;
        RECT 101.125 69.090 101.775 69.120 ;
        RECT 97.995 69.045 98.255 69.090 ;
        RECT 97.160 68.835 97.390 68.980 ;
        RECT 98.800 68.835 99.030 68.980 ;
        RECT 99.730 68.835 99.990 68.910 ;
        RECT 100.735 68.835 100.965 68.980 ;
        RECT 101.935 68.835 102.165 68.980 ;
        RECT 97.160 68.665 102.165 68.835 ;
        RECT 89.995 68.275 91.905 68.380 ;
        RECT 77.465 66.880 78.465 66.910 ;
        RECT 80.995 66.880 81.645 66.910 ;
        RECT 82.235 66.880 82.535 67.135 ;
        RECT 74.265 66.710 75.820 66.775 ;
        RECT 69.870 65.635 70.160 66.710 ;
        RECT 70.755 66.680 71.755 66.710 ;
        RECT 74.285 66.680 74.935 66.710 ;
        RECT 70.735 66.320 70.995 66.365 ;
        RECT 70.735 66.290 71.755 66.320 ;
        RECT 74.285 66.290 74.935 66.320 ;
        RECT 70.735 66.120 74.955 66.290 ;
        RECT 70.735 66.090 71.755 66.120 ;
        RECT 74.285 66.090 74.935 66.120 ;
        RECT 70.735 66.045 70.995 66.090 ;
        RECT 70.320 65.835 70.550 65.980 ;
        RECT 71.960 65.835 72.190 65.980 ;
        RECT 73.895 65.835 74.125 65.980 ;
        RECT 74.695 65.835 74.955 65.910 ;
        RECT 75.095 65.835 75.325 65.980 ;
        RECT 70.320 65.665 75.325 65.835 ;
        RECT 63.155 65.275 65.065 65.380 ;
        RECT 56.450 65.000 56.740 65.210 ;
        RECT 57.335 65.180 58.335 65.210 ;
        RECT 60.865 65.180 61.515 65.210 ;
        RECT 62.110 65.000 62.400 65.210 ;
        RECT 63.160 65.210 65.065 65.275 ;
        RECT 67.555 65.210 69.110 65.380 ;
        RECT 69.865 65.380 70.165 65.635 ;
        RECT 70.320 65.520 70.550 65.665 ;
        RECT 71.960 65.520 72.190 65.665 ;
        RECT 73.895 65.520 74.125 65.665 ;
        RECT 74.695 65.590 74.955 65.665 ;
        RECT 75.095 65.520 75.325 65.665 ;
        RECT 70.755 65.380 71.755 65.410 ;
        RECT 74.285 65.380 74.935 65.410 ;
        RECT 75.530 65.380 75.820 66.710 ;
        RECT 76.580 66.710 78.485 66.880 ;
        RECT 80.975 66.775 82.535 66.880 ;
        RECT 83.290 66.880 83.580 68.210 ;
        RECT 84.175 68.180 85.175 68.210 ;
        RECT 87.705 68.180 88.355 68.210 ;
        RECT 84.995 67.820 85.255 67.865 ;
        RECT 84.175 67.790 85.255 67.820 ;
        RECT 86.310 67.790 86.570 67.865 ;
        RECT 87.705 67.790 88.355 67.820 ;
        RECT 84.155 67.620 88.375 67.790 ;
        RECT 84.175 67.590 85.255 67.620 ;
        RECT 84.995 67.545 85.255 67.590 ;
        RECT 86.310 67.545 86.570 67.620 ;
        RECT 87.705 67.590 88.355 67.620 ;
        RECT 83.740 67.335 83.970 67.480 ;
        RECT 85.380 67.335 85.610 67.480 ;
        RECT 86.280 67.335 86.600 67.380 ;
        RECT 87.315 67.335 87.545 67.480 ;
        RECT 88.515 67.335 88.745 67.480 ;
        RECT 83.740 67.165 88.745 67.335 ;
        RECT 83.740 67.020 83.970 67.165 ;
        RECT 85.380 67.020 85.610 67.165 ;
        RECT 86.280 67.120 86.600 67.165 ;
        RECT 87.315 67.020 87.545 67.165 ;
        RECT 88.515 67.020 88.745 67.165 ;
        RECT 88.950 67.135 89.240 68.210 ;
        RECT 90.000 68.210 91.905 68.275 ;
        RECT 84.175 66.880 85.175 66.910 ;
        RECT 87.705 66.880 88.355 66.910 ;
        RECT 88.945 66.880 89.245 67.135 ;
        RECT 80.975 66.710 82.530 66.775 ;
        RECT 76.580 65.635 76.870 66.710 ;
        RECT 77.465 66.680 78.465 66.710 ;
        RECT 80.995 66.680 81.645 66.710 ;
        RECT 77.465 66.290 78.465 66.320 ;
        RECT 80.995 66.290 81.645 66.320 ;
        RECT 77.445 66.120 81.665 66.290 ;
        RECT 77.465 66.090 78.465 66.120 ;
        RECT 80.995 66.090 81.645 66.120 ;
        RECT 77.030 65.835 77.260 65.980 ;
        RECT 78.670 65.835 78.900 65.980 ;
        RECT 80.605 65.835 80.835 65.980 ;
        RECT 81.805 65.835 82.035 65.980 ;
        RECT 82.240 65.835 82.530 66.710 ;
        RECT 77.030 65.665 82.530 65.835 ;
        RECT 69.865 65.275 71.775 65.380 ;
        RECT 63.160 65.000 63.450 65.210 ;
        RECT 64.045 65.180 65.045 65.210 ;
        RECT 67.575 65.180 68.225 65.210 ;
        RECT 68.820 65.000 69.110 65.210 ;
        RECT 69.870 65.210 71.775 65.275 ;
        RECT 74.265 65.210 75.820 65.380 ;
        RECT 76.575 65.380 76.875 65.635 ;
        RECT 77.030 65.520 77.260 65.665 ;
        RECT 78.670 65.520 78.900 65.665 ;
        RECT 80.605 65.520 80.835 65.665 ;
        RECT 81.805 65.520 82.035 65.665 ;
        RECT 77.465 65.380 78.465 65.410 ;
        RECT 80.995 65.380 81.645 65.410 ;
        RECT 82.240 65.380 82.530 65.665 ;
        RECT 83.290 66.710 85.195 66.880 ;
        RECT 87.685 66.775 89.245 66.880 ;
        RECT 90.000 66.880 90.290 68.210 ;
        RECT 90.885 68.180 91.885 68.210 ;
        RECT 92.130 67.950 92.390 68.270 ;
        RECT 94.395 68.210 95.950 68.380 ;
        RECT 96.705 68.380 97.005 68.635 ;
        RECT 97.160 68.520 97.390 68.665 ;
        RECT 98.800 68.520 99.030 68.665 ;
        RECT 99.730 68.590 99.990 68.665 ;
        RECT 100.735 68.520 100.965 68.665 ;
        RECT 101.935 68.520 102.165 68.665 ;
        RECT 97.595 68.380 98.595 68.410 ;
        RECT 101.125 68.380 101.775 68.410 ;
        RECT 102.370 68.380 102.660 69.710 ;
        RECT 96.705 68.275 98.615 68.380 ;
        RECT 94.415 68.180 95.065 68.210 ;
        RECT 90.885 67.790 91.885 67.820 ;
        RECT 92.175 67.790 92.345 67.950 ;
        RECT 93.020 67.790 93.280 67.865 ;
        RECT 94.415 67.790 95.065 67.820 ;
        RECT 90.865 67.620 95.085 67.790 ;
        RECT 90.885 67.590 91.885 67.620 ;
        RECT 93.020 67.545 93.280 67.620 ;
        RECT 94.415 67.590 95.065 67.620 ;
        RECT 90.450 67.335 90.680 67.480 ;
        RECT 92.090 67.335 92.320 67.480 ;
        RECT 92.990 67.335 93.310 67.380 ;
        RECT 94.025 67.335 94.255 67.480 ;
        RECT 95.225 67.335 95.455 67.480 ;
        RECT 90.450 67.165 95.455 67.335 ;
        RECT 90.450 67.020 90.680 67.165 ;
        RECT 92.090 67.020 92.320 67.165 ;
        RECT 92.990 67.120 93.310 67.165 ;
        RECT 94.025 67.020 94.255 67.165 ;
        RECT 95.225 67.020 95.455 67.165 ;
        RECT 95.660 67.135 95.950 68.210 ;
        RECT 96.710 68.210 98.615 68.275 ;
        RECT 101.105 68.210 102.660 68.380 ;
        RECT 90.885 66.880 91.885 66.910 ;
        RECT 94.415 66.880 95.065 66.910 ;
        RECT 95.655 66.880 95.955 67.135 ;
        RECT 87.685 66.710 89.240 66.775 ;
        RECT 83.290 65.635 83.580 66.710 ;
        RECT 84.175 66.680 85.175 66.710 ;
        RECT 87.705 66.680 88.355 66.710 ;
        RECT 84.155 66.320 84.415 66.365 ;
        RECT 84.155 66.290 85.175 66.320 ;
        RECT 87.705 66.290 88.355 66.320 ;
        RECT 84.155 66.120 88.375 66.290 ;
        RECT 84.155 66.090 85.175 66.120 ;
        RECT 87.705 66.090 88.355 66.120 ;
        RECT 84.155 66.045 84.415 66.090 ;
        RECT 83.740 65.835 83.970 65.980 ;
        RECT 85.380 65.835 85.610 65.980 ;
        RECT 87.315 65.835 87.545 65.980 ;
        RECT 88.115 65.835 88.375 65.910 ;
        RECT 88.515 65.835 88.745 65.980 ;
        RECT 83.740 65.665 88.745 65.835 ;
        RECT 76.575 65.275 78.485 65.380 ;
        RECT 69.870 65.000 70.160 65.210 ;
        RECT 70.755 65.180 71.755 65.210 ;
        RECT 74.285 65.180 74.935 65.210 ;
        RECT 75.530 65.000 75.820 65.210 ;
        RECT 76.580 65.210 78.485 65.275 ;
        RECT 80.975 65.210 82.530 65.380 ;
        RECT 83.285 65.380 83.585 65.635 ;
        RECT 83.740 65.520 83.970 65.665 ;
        RECT 85.380 65.520 85.610 65.665 ;
        RECT 87.315 65.520 87.545 65.665 ;
        RECT 88.115 65.590 88.375 65.665 ;
        RECT 88.515 65.520 88.745 65.665 ;
        RECT 84.175 65.380 85.175 65.410 ;
        RECT 87.705 65.380 88.355 65.410 ;
        RECT 88.950 65.380 89.240 66.710 ;
        RECT 90.000 66.710 91.905 66.880 ;
        RECT 94.395 66.775 95.955 66.880 ;
        RECT 96.710 66.880 97.000 68.210 ;
        RECT 97.595 68.180 98.595 68.210 ;
        RECT 101.125 68.180 101.775 68.210 ;
        RECT 98.415 67.820 98.675 67.865 ;
        RECT 97.595 67.790 98.675 67.820 ;
        RECT 99.730 67.790 99.990 67.865 ;
        RECT 101.125 67.790 101.775 67.820 ;
        RECT 97.575 67.620 101.795 67.790 ;
        RECT 97.595 67.590 98.675 67.620 ;
        RECT 98.415 67.545 98.675 67.590 ;
        RECT 99.730 67.545 99.990 67.620 ;
        RECT 101.125 67.590 101.775 67.620 ;
        RECT 97.160 67.335 97.390 67.480 ;
        RECT 98.800 67.335 99.030 67.480 ;
        RECT 99.700 67.335 100.020 67.380 ;
        RECT 100.735 67.335 100.965 67.480 ;
        RECT 101.935 67.335 102.165 67.480 ;
        RECT 97.160 67.165 102.165 67.335 ;
        RECT 97.160 67.020 97.390 67.165 ;
        RECT 98.800 67.020 99.030 67.165 ;
        RECT 99.700 67.120 100.020 67.165 ;
        RECT 100.735 67.020 100.965 67.165 ;
        RECT 101.935 67.020 102.165 67.165 ;
        RECT 102.370 67.135 102.660 68.210 ;
        RECT 97.595 66.880 98.595 66.910 ;
        RECT 101.125 66.880 101.775 66.910 ;
        RECT 102.365 66.880 102.665 67.135 ;
        RECT 94.395 66.710 95.950 66.775 ;
        RECT 90.000 65.635 90.290 66.710 ;
        RECT 90.885 66.680 91.885 66.710 ;
        RECT 94.415 66.680 95.065 66.710 ;
        RECT 90.885 66.290 91.885 66.320 ;
        RECT 94.415 66.290 95.065 66.320 ;
        RECT 90.865 66.120 95.085 66.290 ;
        RECT 90.885 66.090 91.885 66.120 ;
        RECT 94.415 66.090 95.065 66.120 ;
        RECT 90.450 65.835 90.680 65.980 ;
        RECT 92.090 65.835 92.320 65.980 ;
        RECT 94.025 65.835 94.255 65.980 ;
        RECT 95.225 65.835 95.455 65.980 ;
        RECT 95.660 65.835 95.950 66.710 ;
        RECT 90.450 65.665 95.950 65.835 ;
        RECT 83.285 65.275 85.195 65.380 ;
        RECT 76.580 65.000 76.870 65.210 ;
        RECT 77.465 65.180 78.465 65.210 ;
        RECT 80.995 65.180 81.645 65.210 ;
        RECT 82.240 65.000 82.530 65.210 ;
        RECT 83.290 65.210 85.195 65.275 ;
        RECT 87.685 65.210 89.240 65.380 ;
        RECT 89.995 65.380 90.295 65.635 ;
        RECT 90.450 65.520 90.680 65.665 ;
        RECT 92.090 65.520 92.320 65.665 ;
        RECT 94.025 65.520 94.255 65.665 ;
        RECT 95.225 65.520 95.455 65.665 ;
        RECT 90.885 65.380 91.885 65.410 ;
        RECT 94.415 65.380 95.065 65.410 ;
        RECT 95.660 65.380 95.950 65.665 ;
        RECT 96.710 66.710 98.615 66.880 ;
        RECT 101.105 66.775 102.665 66.880 ;
        RECT 101.105 66.710 102.660 66.775 ;
        RECT 96.710 65.635 97.000 66.710 ;
        RECT 97.595 66.680 98.595 66.710 ;
        RECT 101.125 66.680 101.775 66.710 ;
        RECT 97.575 66.320 97.835 66.365 ;
        RECT 97.575 66.290 98.595 66.320 ;
        RECT 101.125 66.290 101.775 66.320 ;
        RECT 97.575 66.120 101.795 66.290 ;
        RECT 97.575 66.090 98.595 66.120 ;
        RECT 101.125 66.090 101.775 66.120 ;
        RECT 97.575 66.045 97.835 66.090 ;
        RECT 97.160 65.835 97.390 65.980 ;
        RECT 98.800 65.835 99.030 65.980 ;
        RECT 100.735 65.835 100.965 65.980 ;
        RECT 101.535 65.835 101.795 65.910 ;
        RECT 101.935 65.835 102.165 65.980 ;
        RECT 97.160 65.665 102.165 65.835 ;
        RECT 89.995 65.275 91.905 65.380 ;
        RECT 83.290 65.000 83.580 65.210 ;
        RECT 84.175 65.180 85.175 65.210 ;
        RECT 87.705 65.180 88.355 65.210 ;
        RECT 88.950 65.000 89.240 65.210 ;
        RECT 90.000 65.210 91.905 65.275 ;
        RECT 94.395 65.210 95.950 65.380 ;
        RECT 96.705 65.380 97.005 65.635 ;
        RECT 97.160 65.520 97.390 65.665 ;
        RECT 98.800 65.520 99.030 65.665 ;
        RECT 100.735 65.520 100.965 65.665 ;
        RECT 101.535 65.590 101.795 65.665 ;
        RECT 101.935 65.520 102.165 65.665 ;
        RECT 97.595 65.380 98.595 65.410 ;
        RECT 101.125 65.380 101.775 65.410 ;
        RECT 102.370 65.380 102.660 66.710 ;
        RECT 96.705 65.275 98.615 65.380 ;
        RECT 90.000 65.000 90.290 65.210 ;
        RECT 90.885 65.180 91.885 65.210 ;
        RECT 94.415 65.180 95.065 65.210 ;
        RECT 95.660 65.000 95.950 65.210 ;
        RECT 96.710 65.210 98.615 65.275 ;
        RECT 101.105 65.210 102.660 65.380 ;
        RECT 96.710 65.000 97.000 65.210 ;
        RECT 97.595 65.180 98.595 65.210 ;
        RECT 101.125 65.180 101.775 65.210 ;
        RECT 102.370 65.000 102.660 65.210 ;
        RECT 47.855 64.830 48.115 64.905 ;
        RECT 92.600 64.830 92.860 64.905 ;
        RECT 47.855 64.660 92.860 64.830 ;
        RECT 47.855 64.585 48.115 64.660 ;
        RECT 92.600 64.585 92.860 64.660 ;
        RECT 61.275 64.445 61.535 64.520 ;
        RECT 89.535 64.445 89.795 64.520 ;
        RECT 61.275 64.275 89.795 64.445 ;
        RECT 61.275 64.200 61.535 64.275 ;
        RECT 89.535 64.200 89.795 64.275 ;
        RECT 74.695 64.060 74.955 64.135 ;
        RECT 99.310 64.060 99.570 64.135 ;
        RECT 74.695 63.890 99.570 64.060 ;
        RECT 74.695 63.815 74.955 63.890 ;
        RECT 99.310 63.815 99.570 63.890 ;
        RECT 39.340 63.675 39.600 63.750 ;
        RECT 52.760 63.675 53.020 63.750 ;
        RECT 66.150 63.675 66.470 63.720 ;
        RECT 79.600 63.675 79.860 63.750 ;
        RECT 39.340 63.505 79.860 63.675 ;
        RECT 39.340 63.430 39.600 63.505 ;
        RECT 52.760 63.430 53.020 63.505 ;
        RECT 66.150 63.460 66.470 63.505 ;
        RECT 79.600 63.430 79.860 63.505 ;
        RECT 88.115 63.675 88.375 63.750 ;
        RECT 96.245 63.675 96.505 63.750 ;
        RECT 88.115 63.505 96.505 63.675 ;
        RECT 88.115 63.430 88.375 63.505 ;
        RECT 96.245 63.430 96.505 63.505 ;
        RECT 46.050 63.290 46.310 63.365 ;
        RECT 59.470 63.290 59.730 63.365 ;
        RECT 72.890 63.290 73.150 63.365 ;
        RECT 86.310 63.290 86.570 63.365 ;
        RECT 46.050 63.120 86.570 63.290 ;
        RECT 46.050 63.045 46.310 63.120 ;
        RECT 59.470 63.045 59.730 63.120 ;
        RECT 72.890 63.045 73.150 63.120 ;
        RECT 86.310 63.045 86.570 63.120 ;
        RECT 0.000 0.000 1.000 1.000 ;
        RECT 144.360 0.000 145.360 1.000 ;
      LAYER met2 ;
        RECT 17.600 198.395 18.100 207.880 ;
        RECT 18.350 201.920 18.850 207.880 ;
        RECT 19.655 203.150 19.935 203.205 ;
        RECT 21.155 203.150 21.435 203.205 ;
        RECT 22.655 203.150 22.935 203.205 ;
        RECT 24.155 203.150 24.435 203.205 ;
        RECT 25.655 203.150 25.935 203.205 ;
        RECT 27.155 203.150 27.435 203.205 ;
        RECT 28.655 203.150 28.935 203.205 ;
        RECT 30.155 203.150 30.435 203.205 ;
        RECT 19.635 202.890 19.955 203.150 ;
        RECT 21.135 202.890 21.455 203.150 ;
        RECT 22.635 202.890 22.955 203.150 ;
        RECT 24.135 202.890 24.455 203.150 ;
        RECT 25.635 202.890 25.955 203.150 ;
        RECT 27.135 202.890 27.455 203.150 ;
        RECT 28.635 202.890 28.955 203.150 ;
        RECT 30.135 202.890 30.455 203.150 ;
        RECT 19.655 202.835 19.935 202.890 ;
        RECT 21.155 202.835 21.435 202.890 ;
        RECT 22.655 202.835 22.935 202.890 ;
        RECT 24.155 202.835 24.435 202.890 ;
        RECT 25.655 202.835 25.935 202.890 ;
        RECT 27.155 202.835 27.435 202.890 ;
        RECT 28.655 202.835 28.935 202.890 ;
        RECT 30.155 202.835 30.435 202.890 ;
        RECT 30.830 201.920 31.330 207.880 ;
        RECT 18.350 201.420 19.350 201.920 ;
        RECT 18.850 200.395 19.350 201.420 ;
        RECT 30.330 201.420 31.330 201.920 ;
        RECT 30.330 200.395 30.830 201.420 ;
        RECT 18.580 199.445 19.620 200.395 ;
        RECT 30.060 199.445 31.100 200.395 ;
        RECT 31.580 198.395 32.080 207.880 ;
        RECT 39.680 198.395 40.180 207.880 ;
        RECT 40.430 201.920 40.930 207.880 ;
        RECT 41.735 203.150 42.015 203.205 ;
        RECT 43.235 203.150 43.515 203.205 ;
        RECT 44.735 203.150 45.015 203.205 ;
        RECT 46.235 203.150 46.515 203.205 ;
        RECT 47.735 203.150 48.015 203.205 ;
        RECT 49.235 203.150 49.515 203.205 ;
        RECT 50.735 203.150 51.015 203.205 ;
        RECT 52.235 203.150 52.515 203.205 ;
        RECT 41.715 202.890 42.035 203.150 ;
        RECT 43.215 202.890 43.535 203.150 ;
        RECT 44.715 202.890 45.035 203.150 ;
        RECT 46.215 202.890 46.535 203.150 ;
        RECT 47.715 202.890 48.035 203.150 ;
        RECT 49.215 202.890 49.535 203.150 ;
        RECT 50.715 202.890 51.035 203.150 ;
        RECT 52.215 202.890 52.535 203.150 ;
        RECT 41.735 202.835 42.015 202.890 ;
        RECT 43.235 202.835 43.515 202.890 ;
        RECT 44.735 202.835 45.015 202.890 ;
        RECT 46.235 202.835 46.515 202.890 ;
        RECT 47.735 202.835 48.015 202.890 ;
        RECT 49.235 202.835 49.515 202.890 ;
        RECT 50.735 202.835 51.015 202.890 ;
        RECT 52.235 202.835 52.515 202.890 ;
        RECT 52.910 201.920 53.410 207.880 ;
        RECT 40.430 201.420 41.430 201.920 ;
        RECT 40.930 200.395 41.430 201.420 ;
        RECT 52.410 201.420 53.410 201.920 ;
        RECT 52.410 200.395 52.910 201.420 ;
        RECT 40.660 199.445 41.700 200.395 ;
        RECT 52.140 199.445 53.180 200.395 ;
        RECT 53.660 198.395 54.160 207.880 ;
        RECT 61.760 198.395 62.260 207.880 ;
        RECT 62.510 201.920 63.010 207.880 ;
        RECT 63.815 203.150 64.095 203.205 ;
        RECT 65.315 203.150 65.595 203.205 ;
        RECT 66.815 203.150 67.095 203.205 ;
        RECT 68.315 203.150 68.595 203.205 ;
        RECT 69.815 203.150 70.095 203.205 ;
        RECT 71.315 203.150 71.595 203.205 ;
        RECT 72.815 203.150 73.095 203.205 ;
        RECT 74.315 203.150 74.595 203.205 ;
        RECT 63.795 202.890 64.115 203.150 ;
        RECT 65.295 202.890 65.615 203.150 ;
        RECT 66.795 202.890 67.115 203.150 ;
        RECT 68.295 202.890 68.615 203.150 ;
        RECT 69.795 202.890 70.115 203.150 ;
        RECT 71.295 202.890 71.615 203.150 ;
        RECT 72.795 202.890 73.115 203.150 ;
        RECT 74.295 202.890 74.615 203.150 ;
        RECT 63.815 202.835 64.095 202.890 ;
        RECT 65.315 202.835 65.595 202.890 ;
        RECT 66.815 202.835 67.095 202.890 ;
        RECT 68.315 202.835 68.595 202.890 ;
        RECT 69.815 202.835 70.095 202.890 ;
        RECT 71.315 202.835 71.595 202.890 ;
        RECT 72.815 202.835 73.095 202.890 ;
        RECT 74.315 202.835 74.595 202.890 ;
        RECT 74.990 201.920 75.490 207.880 ;
        RECT 62.510 201.420 63.510 201.920 ;
        RECT 63.010 200.395 63.510 201.420 ;
        RECT 74.490 201.420 75.490 201.920 ;
        RECT 74.490 200.395 74.990 201.420 ;
        RECT 62.740 199.445 63.780 200.395 ;
        RECT 74.220 199.445 75.260 200.395 ;
        RECT 75.740 198.395 76.240 207.880 ;
        RECT 105.620 202.420 106.120 207.880 ;
        RECT 106.370 204.420 106.870 207.880 ;
        RECT 107.735 207.090 108.015 207.145 ;
        RECT 109.235 207.090 109.515 207.145 ;
        RECT 110.735 207.090 111.015 207.145 ;
        RECT 112.235 207.090 112.515 207.145 ;
        RECT 113.735 207.090 114.015 207.145 ;
        RECT 115.235 207.090 115.515 207.145 ;
        RECT 116.735 207.090 117.015 207.145 ;
        RECT 118.235 207.090 118.515 207.145 ;
        RECT 107.715 206.830 108.035 207.090 ;
        RECT 109.215 206.830 109.535 207.090 ;
        RECT 110.715 206.830 111.035 207.090 ;
        RECT 112.215 206.830 112.535 207.090 ;
        RECT 113.715 206.830 114.035 207.090 ;
        RECT 115.215 206.830 115.535 207.090 ;
        RECT 116.715 206.830 117.035 207.090 ;
        RECT 118.215 206.830 118.535 207.090 ;
        RECT 107.735 206.775 108.015 206.830 ;
        RECT 109.235 206.775 109.515 206.830 ;
        RECT 110.735 206.775 111.015 206.830 ;
        RECT 112.235 206.775 112.515 206.830 ;
        RECT 113.735 206.775 114.015 206.830 ;
        RECT 115.235 206.775 115.515 206.830 ;
        RECT 116.735 206.775 117.015 206.830 ;
        RECT 118.235 206.775 118.515 206.830 ;
        RECT 119.445 204.420 119.945 207.880 ;
        RECT 106.370 203.420 107.415 204.420 ;
        RECT 118.900 203.420 119.945 204.420 ;
        RECT 105.120 201.420 106.165 202.420 ;
        RECT 106.370 201.605 106.870 203.420 ;
        RECT 108.200 202.470 108.460 202.790 ;
        RECT 109.700 202.470 109.960 202.790 ;
        RECT 111.200 202.470 111.460 202.790 ;
        RECT 112.700 202.470 112.960 202.790 ;
        RECT 114.200 202.470 114.460 202.790 ;
        RECT 115.700 202.470 115.960 202.790 ;
        RECT 117.200 202.470 117.460 202.790 ;
        RECT 118.700 202.470 118.960 202.790 ;
        RECT 107.745 202.050 108.005 202.370 ;
        RECT 17.330 197.445 18.370 198.395 ;
        RECT 31.310 197.445 32.350 198.395 ;
        RECT 39.410 197.445 40.450 198.395 ;
        RECT 53.390 197.445 54.430 198.395 ;
        RECT 61.490 197.445 62.530 198.395 ;
        RECT 75.470 197.445 76.510 198.395 ;
        RECT 105.620 188.000 106.120 201.420 ;
        RECT 106.370 200.420 106.870 200.870 ;
        RECT 106.370 199.420 107.415 200.420 ;
        RECT 106.370 188.000 106.870 199.420 ;
        RECT 107.260 198.110 107.580 198.155 ;
        RECT 107.790 198.110 107.960 202.050 ;
        RECT 107.260 197.940 107.960 198.110 ;
        RECT 107.260 197.895 107.580 197.940 ;
        RECT 108.245 197.645 108.415 202.470 ;
        RECT 109.245 202.050 109.505 202.370 ;
        RECT 108.760 198.110 109.080 198.155 ;
        RECT 109.290 198.110 109.460 202.050 ;
        RECT 108.760 197.940 109.460 198.110 ;
        RECT 108.760 197.895 109.080 197.940 ;
        RECT 109.745 197.645 109.915 202.470 ;
        RECT 110.745 202.050 111.005 202.370 ;
        RECT 110.260 198.110 110.580 198.155 ;
        RECT 110.790 198.110 110.960 202.050 ;
        RECT 110.260 197.940 110.960 198.110 ;
        RECT 110.260 197.895 110.580 197.940 ;
        RECT 111.245 197.645 111.415 202.470 ;
        RECT 112.245 202.050 112.505 202.370 ;
        RECT 111.760 198.110 112.080 198.155 ;
        RECT 112.290 198.110 112.460 202.050 ;
        RECT 111.760 197.940 112.460 198.110 ;
        RECT 111.760 197.895 112.080 197.940 ;
        RECT 112.745 197.645 112.915 202.470 ;
        RECT 113.745 202.050 114.005 202.370 ;
        RECT 113.260 198.110 113.580 198.155 ;
        RECT 113.790 198.110 113.960 202.050 ;
        RECT 113.260 197.940 113.960 198.110 ;
        RECT 113.260 197.895 113.580 197.940 ;
        RECT 114.245 197.645 114.415 202.470 ;
        RECT 115.245 202.050 115.505 202.370 ;
        RECT 114.760 198.110 115.080 198.155 ;
        RECT 115.290 198.110 115.460 202.050 ;
        RECT 114.760 197.940 115.460 198.110 ;
        RECT 114.760 197.895 115.080 197.940 ;
        RECT 115.745 197.645 115.915 202.470 ;
        RECT 116.745 202.050 117.005 202.370 ;
        RECT 116.260 198.110 116.580 198.155 ;
        RECT 116.790 198.110 116.960 202.050 ;
        RECT 116.260 197.940 116.960 198.110 ;
        RECT 116.260 197.895 116.580 197.940 ;
        RECT 117.245 197.645 117.415 202.470 ;
        RECT 118.245 202.050 118.505 202.370 ;
        RECT 117.760 198.110 118.080 198.155 ;
        RECT 118.290 198.110 118.460 202.050 ;
        RECT 117.760 197.940 118.460 198.110 ;
        RECT 117.760 197.895 118.080 197.940 ;
        RECT 118.745 197.645 118.915 202.470 ;
        RECT 119.445 201.605 119.945 203.420 ;
        RECT 120.195 202.420 120.695 207.880 ;
        RECT 120.150 201.420 121.195 202.420 ;
        RECT 107.335 197.475 108.415 197.645 ;
        RECT 108.835 197.475 109.915 197.645 ;
        RECT 110.335 197.475 111.415 197.645 ;
        RECT 111.835 197.475 112.915 197.645 ;
        RECT 113.335 197.475 114.415 197.645 ;
        RECT 114.835 197.475 115.915 197.645 ;
        RECT 116.335 197.475 117.415 197.645 ;
        RECT 117.835 197.475 118.915 197.645 ;
        RECT 107.335 190.975 107.505 197.475 ;
        RECT 107.745 196.945 108.005 197.265 ;
        RECT 107.790 193.165 107.960 196.945 ;
        RECT 108.170 195.790 108.490 196.050 ;
        RECT 108.245 193.725 108.415 195.790 ;
        RECT 108.245 193.480 108.555 193.725 ;
        RECT 108.295 193.405 108.555 193.480 ;
        RECT 108.200 193.165 108.460 193.240 ;
        RECT 107.790 192.995 108.460 193.165 ;
        RECT 108.200 192.920 108.460 192.995 ;
        RECT 108.835 190.975 109.005 197.475 ;
        RECT 109.245 196.945 109.505 197.265 ;
        RECT 109.290 193.165 109.460 196.945 ;
        RECT 109.670 195.790 109.990 196.050 ;
        RECT 109.745 193.725 109.915 195.790 ;
        RECT 109.745 193.480 110.055 193.725 ;
        RECT 109.795 193.405 110.055 193.480 ;
        RECT 109.700 193.165 109.960 193.240 ;
        RECT 109.290 192.995 109.960 193.165 ;
        RECT 109.700 192.920 109.960 192.995 ;
        RECT 110.335 190.975 110.505 197.475 ;
        RECT 110.745 196.945 111.005 197.265 ;
        RECT 110.790 193.165 110.960 196.945 ;
        RECT 111.170 195.790 111.490 196.050 ;
        RECT 111.245 193.725 111.415 195.790 ;
        RECT 111.245 193.480 111.555 193.725 ;
        RECT 111.295 193.405 111.555 193.480 ;
        RECT 111.200 193.165 111.460 193.240 ;
        RECT 110.790 192.995 111.460 193.165 ;
        RECT 111.200 192.920 111.460 192.995 ;
        RECT 111.835 190.975 112.005 197.475 ;
        RECT 112.245 196.945 112.505 197.265 ;
        RECT 112.290 193.165 112.460 196.945 ;
        RECT 112.670 195.790 112.990 196.050 ;
        RECT 112.745 193.725 112.915 195.790 ;
        RECT 112.745 193.480 113.055 193.725 ;
        RECT 112.795 193.405 113.055 193.480 ;
        RECT 112.700 193.165 112.960 193.240 ;
        RECT 112.290 192.995 112.960 193.165 ;
        RECT 112.700 192.920 112.960 192.995 ;
        RECT 113.335 190.975 113.505 197.475 ;
        RECT 113.745 196.945 114.005 197.265 ;
        RECT 113.790 193.165 113.960 196.945 ;
        RECT 114.170 195.790 114.490 196.050 ;
        RECT 114.245 193.725 114.415 195.790 ;
        RECT 114.245 193.480 114.555 193.725 ;
        RECT 114.295 193.405 114.555 193.480 ;
        RECT 114.200 193.165 114.460 193.240 ;
        RECT 113.790 192.995 114.460 193.165 ;
        RECT 114.200 192.920 114.460 192.995 ;
        RECT 114.835 190.975 115.005 197.475 ;
        RECT 115.245 196.945 115.505 197.265 ;
        RECT 115.290 193.165 115.460 196.945 ;
        RECT 115.670 195.790 115.990 196.050 ;
        RECT 115.745 193.725 115.915 195.790 ;
        RECT 115.745 193.480 116.055 193.725 ;
        RECT 115.795 193.405 116.055 193.480 ;
        RECT 115.700 193.165 115.960 193.240 ;
        RECT 115.290 192.995 115.960 193.165 ;
        RECT 115.700 192.920 115.960 192.995 ;
        RECT 116.335 190.975 116.505 197.475 ;
        RECT 116.745 196.945 117.005 197.265 ;
        RECT 116.790 193.165 116.960 196.945 ;
        RECT 117.170 195.790 117.490 196.050 ;
        RECT 117.245 193.725 117.415 195.790 ;
        RECT 117.245 193.480 117.555 193.725 ;
        RECT 117.295 193.405 117.555 193.480 ;
        RECT 117.200 193.165 117.460 193.240 ;
        RECT 116.790 192.995 117.460 193.165 ;
        RECT 117.200 192.920 117.460 192.995 ;
        RECT 117.835 190.975 118.005 197.475 ;
        RECT 118.245 196.945 118.505 197.265 ;
        RECT 118.290 193.165 118.460 196.945 ;
        RECT 118.670 195.790 118.990 196.050 ;
        RECT 118.745 193.725 118.915 195.790 ;
        RECT 118.745 193.480 119.055 193.725 ;
        RECT 118.795 193.405 119.055 193.480 ;
        RECT 118.700 193.165 118.960 193.240 ;
        RECT 118.290 192.995 118.960 193.165 ;
        RECT 118.700 192.920 118.960 192.995 ;
        RECT 119.445 192.420 119.945 200.870 ;
        RECT 118.900 191.420 119.945 192.420 ;
        RECT 107.335 190.805 107.960 190.975 ;
        RECT 108.835 190.805 109.460 190.975 ;
        RECT 110.335 190.805 110.960 190.975 ;
        RECT 111.835 190.805 112.460 190.975 ;
        RECT 113.335 190.805 113.960 190.975 ;
        RECT 114.835 190.805 115.460 190.975 ;
        RECT 116.335 190.805 116.960 190.975 ;
        RECT 117.835 190.805 118.460 190.975 ;
        RECT 107.790 190.120 107.960 190.805 ;
        RECT 109.290 190.120 109.460 190.805 ;
        RECT 110.790 190.120 110.960 190.805 ;
        RECT 112.290 190.120 112.460 190.805 ;
        RECT 113.790 190.120 113.960 190.805 ;
        RECT 115.290 190.120 115.460 190.805 ;
        RECT 116.790 190.120 116.960 190.805 ;
        RECT 118.290 190.120 118.460 190.805 ;
        RECT 107.715 189.860 108.035 190.120 ;
        RECT 109.215 189.860 109.535 190.120 ;
        RECT 110.715 189.860 111.035 190.120 ;
        RECT 112.215 189.860 112.535 190.120 ;
        RECT 113.715 189.860 114.035 190.120 ;
        RECT 115.215 189.860 115.535 190.120 ;
        RECT 116.715 189.860 117.035 190.120 ;
        RECT 118.215 189.860 118.535 190.120 ;
        RECT 108.190 189.310 108.470 189.365 ;
        RECT 109.690 189.310 109.970 189.365 ;
        RECT 111.190 189.310 111.470 189.365 ;
        RECT 112.690 189.310 112.970 189.365 ;
        RECT 114.190 189.310 114.470 189.365 ;
        RECT 115.690 189.310 115.970 189.365 ;
        RECT 117.190 189.310 117.470 189.365 ;
        RECT 118.690 189.310 118.970 189.365 ;
        RECT 108.170 189.050 108.490 189.310 ;
        RECT 109.670 189.050 109.990 189.310 ;
        RECT 111.170 189.050 111.490 189.310 ;
        RECT 112.670 189.050 112.990 189.310 ;
        RECT 114.170 189.050 114.490 189.310 ;
        RECT 115.670 189.050 115.990 189.310 ;
        RECT 117.170 189.050 117.490 189.310 ;
        RECT 118.670 189.050 118.990 189.310 ;
        RECT 108.190 188.995 108.470 189.050 ;
        RECT 109.690 188.995 109.970 189.050 ;
        RECT 111.190 188.995 111.470 189.050 ;
        RECT 112.690 188.995 112.970 189.050 ;
        RECT 114.190 188.995 114.470 189.050 ;
        RECT 115.690 188.995 115.970 189.050 ;
        RECT 117.190 188.995 117.470 189.050 ;
        RECT 118.690 188.995 118.970 189.050 ;
        RECT 119.445 188.000 119.945 191.420 ;
        RECT 120.195 188.000 120.695 201.420 ;
        RECT 113.485 165.855 113.765 165.955 ;
        RECT 54.435 165.685 113.765 165.855 ;
        RECT 34.615 163.070 34.975 163.370 ;
        RECT 32.775 159.670 33.815 160.620 ;
        RECT 33.145 157.710 33.445 159.670 ;
        RECT 34.645 158.620 34.945 163.070 ;
        RECT 54.435 162.915 54.605 165.685 ;
        RECT 113.485 165.585 113.765 165.685 ;
        RECT 112.855 165.445 113.135 165.545 ;
        RECT 67.915 165.275 113.135 165.445 ;
        RECT 67.915 162.915 68.085 165.275 ;
        RECT 112.855 165.175 113.135 165.275 ;
        RECT 114.745 165.035 115.025 165.135 ;
        RECT 81.395 164.865 115.025 165.035 ;
        RECT 81.395 162.915 81.565 164.865 ;
        RECT 114.745 164.765 115.025 164.865 ;
        RECT 112.225 164.625 112.505 164.725 ;
        RECT 93.375 164.455 112.505 164.625 ;
        RECT 93.375 162.945 93.545 164.455 ;
        RECT 112.225 164.355 112.505 164.455 ;
        RECT 114.115 164.215 114.395 164.315 ;
        RECT 94.875 164.045 114.395 164.215 ;
        RECT 54.390 162.595 54.650 162.915 ;
        RECT 67.870 162.595 68.130 162.915 ;
        RECT 81.350 162.595 81.610 162.915 ;
        RECT 93.330 162.625 93.590 162.945 ;
        RECT 94.875 162.915 95.045 164.045 ;
        RECT 114.115 163.945 114.395 164.045 ;
        RECT 103.655 163.070 104.015 163.370 ;
        RECT 94.830 162.595 95.090 162.915 ;
        RECT 46.890 162.030 47.150 162.105 ;
        RECT 52.435 162.030 52.695 162.105 ;
        RECT 46.890 161.860 52.695 162.030 ;
        RECT 46.890 161.785 47.150 161.860 ;
        RECT 52.435 161.785 52.695 161.860 ;
        RECT 60.370 162.030 60.630 162.105 ;
        RECT 65.915 162.030 66.175 162.105 ;
        RECT 60.370 161.860 66.175 162.030 ;
        RECT 60.370 161.785 60.630 161.860 ;
        RECT 65.915 161.785 66.175 161.860 ;
        RECT 73.850 162.030 74.110 162.105 ;
        RECT 79.395 162.030 79.655 162.105 ;
        RECT 73.850 161.860 79.655 162.030 ;
        RECT 73.850 161.785 74.110 161.860 ;
        RECT 79.395 161.785 79.655 161.860 ;
        RECT 87.330 162.030 87.590 162.105 ;
        RECT 92.875 162.030 93.135 162.105 ;
        RECT 87.330 161.860 93.135 162.030 ;
        RECT 87.330 161.785 87.590 161.860 ;
        RECT 92.875 161.785 93.135 161.860 ;
        RECT 48.390 161.110 48.650 161.185 ;
        RECT 53.935 161.110 54.195 161.185 ;
        RECT 48.390 160.940 54.195 161.110 ;
        RECT 48.390 160.865 48.650 160.940 ;
        RECT 53.935 160.865 54.195 160.940 ;
        RECT 61.870 161.110 62.130 161.185 ;
        RECT 67.415 161.110 67.675 161.185 ;
        RECT 61.870 160.940 67.675 161.110 ;
        RECT 61.870 160.865 62.130 160.940 ;
        RECT 67.415 160.865 67.675 160.940 ;
        RECT 75.350 161.110 75.610 161.185 ;
        RECT 80.895 161.110 81.155 161.185 ;
        RECT 75.350 160.940 81.155 161.110 ;
        RECT 75.350 160.865 75.610 160.940 ;
        RECT 80.895 160.865 81.155 160.940 ;
        RECT 88.830 161.110 89.090 161.185 ;
        RECT 94.375 161.110 94.635 161.185 ;
        RECT 88.830 160.940 94.635 161.110 ;
        RECT 88.830 160.865 89.090 160.940 ;
        RECT 94.375 160.865 94.635 160.940 ;
        RECT 43.435 160.650 43.695 160.725 ;
        RECT 44.935 160.650 45.195 160.725 ;
        RECT 43.435 160.480 45.195 160.650 ;
        RECT 43.435 160.405 43.695 160.480 ;
        RECT 44.935 160.405 45.195 160.480 ;
        RECT 46.435 160.650 46.695 160.725 ;
        RECT 47.935 160.650 48.195 160.725 ;
        RECT 46.435 160.480 48.195 160.650 ;
        RECT 46.435 160.405 46.695 160.480 ;
        RECT 47.935 160.405 48.195 160.480 ;
        RECT 49.435 160.650 49.695 160.725 ;
        RECT 50.935 160.650 51.195 160.725 ;
        RECT 49.435 160.480 51.195 160.650 ;
        RECT 49.435 160.405 49.695 160.480 ;
        RECT 50.935 160.405 51.195 160.480 ;
        RECT 56.915 160.650 57.175 160.725 ;
        RECT 58.415 160.650 58.675 160.725 ;
        RECT 56.915 160.480 58.675 160.650 ;
        RECT 56.915 160.405 57.175 160.480 ;
        RECT 58.415 160.405 58.675 160.480 ;
        RECT 59.915 160.650 60.175 160.725 ;
        RECT 61.415 160.650 61.675 160.725 ;
        RECT 59.915 160.480 61.675 160.650 ;
        RECT 59.915 160.405 60.175 160.480 ;
        RECT 61.415 160.405 61.675 160.480 ;
        RECT 62.915 160.650 63.175 160.725 ;
        RECT 64.415 160.650 64.675 160.725 ;
        RECT 62.915 160.480 64.675 160.650 ;
        RECT 62.915 160.405 63.175 160.480 ;
        RECT 64.415 160.405 64.675 160.480 ;
        RECT 70.395 160.650 70.655 160.725 ;
        RECT 71.895 160.650 72.155 160.725 ;
        RECT 70.395 160.480 72.155 160.650 ;
        RECT 70.395 160.405 70.655 160.480 ;
        RECT 71.895 160.405 72.155 160.480 ;
        RECT 73.395 160.650 73.655 160.725 ;
        RECT 74.895 160.650 75.155 160.725 ;
        RECT 73.395 160.480 75.155 160.650 ;
        RECT 73.395 160.405 73.655 160.480 ;
        RECT 74.895 160.405 75.155 160.480 ;
        RECT 76.395 160.650 76.655 160.725 ;
        RECT 77.895 160.650 78.155 160.725 ;
        RECT 76.395 160.480 78.155 160.650 ;
        RECT 76.395 160.405 76.655 160.480 ;
        RECT 77.895 160.405 78.155 160.480 ;
        RECT 83.875 160.650 84.135 160.725 ;
        RECT 85.375 160.650 85.635 160.725 ;
        RECT 83.875 160.480 85.635 160.650 ;
        RECT 83.875 160.405 84.135 160.480 ;
        RECT 85.375 160.405 85.635 160.480 ;
        RECT 86.875 160.650 87.135 160.725 ;
        RECT 88.375 160.650 88.635 160.725 ;
        RECT 86.875 160.480 88.635 160.650 ;
        RECT 86.875 160.405 87.135 160.480 ;
        RECT 88.375 160.405 88.635 160.480 ;
        RECT 89.875 160.650 90.135 160.725 ;
        RECT 91.375 160.650 91.635 160.725 ;
        RECT 89.875 160.480 91.635 160.650 ;
        RECT 89.875 160.405 90.135 160.480 ;
        RECT 91.375 160.405 91.635 160.480 ;
        RECT 33.115 157.410 33.475 157.710 ;
        RECT 34.275 157.670 35.315 158.620 ;
        RECT 33.145 154.010 33.445 157.410 ;
        RECT 33.110 153.730 33.480 154.010 ;
        RECT 33.145 151.010 33.445 153.730 ;
        RECT 34.645 152.510 34.945 157.670 ;
        RECT 43.480 156.590 43.650 160.405 ;
        RECT 43.890 160.190 44.150 160.265 ;
        RECT 46.435 160.190 46.695 160.265 ;
        RECT 43.890 160.020 46.695 160.190 ;
        RECT 43.890 159.945 44.150 160.020 ;
        RECT 46.435 159.945 46.695 160.020 ;
        RECT 49.890 160.190 50.150 160.265 ;
        RECT 52.890 160.190 53.150 160.265 ;
        RECT 49.890 160.020 53.150 160.190 ;
        RECT 49.890 159.945 50.150 160.020 ;
        RECT 52.890 159.945 53.150 160.020 ;
        RECT 45.390 159.270 45.650 159.345 ;
        RECT 49.435 159.270 49.695 159.345 ;
        RECT 45.390 159.100 49.695 159.270 ;
        RECT 45.390 159.025 45.650 159.100 ;
        RECT 49.435 159.025 49.695 159.100 ;
        RECT 49.935 156.990 50.105 159.945 ;
        RECT 51.390 159.270 51.650 159.345 ;
        RECT 54.390 159.270 54.650 159.345 ;
        RECT 51.390 159.100 54.650 159.270 ;
        RECT 51.390 159.025 51.650 159.100 ;
        RECT 54.390 159.025 54.650 159.100 ;
        RECT 49.860 156.730 50.180 156.990 ;
        RECT 56.960 156.930 57.130 160.405 ;
        RECT 57.370 160.190 57.630 160.265 ;
        RECT 59.915 160.190 60.175 160.265 ;
        RECT 57.370 160.020 60.175 160.190 ;
        RECT 57.370 159.945 57.630 160.020 ;
        RECT 59.915 159.945 60.175 160.020 ;
        RECT 63.370 160.190 63.630 160.265 ;
        RECT 66.370 160.190 66.630 160.265 ;
        RECT 63.370 160.020 66.630 160.190 ;
        RECT 63.370 159.945 63.630 160.020 ;
        RECT 66.370 159.945 66.630 160.020 ;
        RECT 58.870 159.270 59.130 159.345 ;
        RECT 62.915 159.270 63.175 159.345 ;
        RECT 58.870 159.100 63.175 159.270 ;
        RECT 58.870 159.025 59.130 159.100 ;
        RECT 62.915 159.025 63.175 159.100 ;
        RECT 63.415 157.315 63.585 159.945 ;
        RECT 64.870 159.270 65.130 159.345 ;
        RECT 67.870 159.270 68.130 159.345 ;
        RECT 64.870 159.100 68.130 159.270 ;
        RECT 64.870 159.025 65.130 159.100 ;
        RECT 67.870 159.025 68.130 159.100 ;
        RECT 58.220 157.145 63.585 157.315 ;
        RECT 58.220 156.990 58.390 157.145 ;
        RECT 51.895 156.760 57.130 156.930 ;
        RECT 51.895 156.590 52.065 156.760 ;
        RECT 58.145 156.730 58.465 156.990 ;
        RECT 70.440 156.930 70.610 160.405 ;
        RECT 70.850 160.190 71.110 160.265 ;
        RECT 73.395 160.190 73.655 160.265 ;
        RECT 70.850 160.020 73.655 160.190 ;
        RECT 70.850 159.945 71.110 160.020 ;
        RECT 73.395 159.945 73.655 160.020 ;
        RECT 76.850 160.190 77.110 160.265 ;
        RECT 79.850 160.190 80.110 160.265 ;
        RECT 76.850 160.020 80.110 160.190 ;
        RECT 76.850 159.945 77.110 160.020 ;
        RECT 79.850 159.945 80.110 160.020 ;
        RECT 72.350 159.270 72.610 159.345 ;
        RECT 76.395 159.270 76.655 159.345 ;
        RECT 72.350 159.100 76.655 159.270 ;
        RECT 72.350 159.025 72.610 159.100 ;
        RECT 76.395 159.025 76.655 159.100 ;
        RECT 76.895 157.020 77.065 159.945 ;
        RECT 78.350 159.270 78.610 159.345 ;
        RECT 81.350 159.270 81.610 159.345 ;
        RECT 78.350 159.100 81.610 159.270 ;
        RECT 78.350 159.025 78.610 159.100 ;
        RECT 81.350 159.025 81.610 159.100 ;
        RECT 58.605 156.760 70.610 156.930 ;
        RECT 76.820 156.760 77.140 157.020 ;
        RECT 58.605 156.590 58.775 156.760 ;
        RECT 83.920 156.590 84.090 160.405 ;
        RECT 84.330 160.190 84.590 160.265 ;
        RECT 86.875 160.190 87.135 160.265 ;
        RECT 84.330 160.020 87.135 160.190 ;
        RECT 84.330 159.945 84.590 160.020 ;
        RECT 86.875 159.945 87.135 160.020 ;
        RECT 90.330 160.190 90.590 160.265 ;
        RECT 93.330 160.190 93.590 160.265 ;
        RECT 90.330 160.020 93.590 160.190 ;
        RECT 90.330 159.945 90.590 160.020 ;
        RECT 93.330 159.945 93.590 160.020 ;
        RECT 85.830 159.270 86.090 159.345 ;
        RECT 89.875 159.270 90.135 159.345 ;
        RECT 85.830 159.100 90.135 159.270 ;
        RECT 85.830 159.025 86.090 159.100 ;
        RECT 89.875 159.025 90.135 159.100 ;
        RECT 90.375 156.975 90.545 159.945 ;
        RECT 91.830 159.270 92.090 159.345 ;
        RECT 94.830 159.270 95.090 159.345 ;
        RECT 91.830 159.100 95.090 159.270 ;
        RECT 91.830 159.025 92.090 159.100 ;
        RECT 94.830 159.025 95.090 159.100 ;
        RECT 103.685 158.620 103.985 163.070 ;
        RECT 104.815 159.670 105.855 160.620 ;
        RECT 103.320 157.670 104.360 158.620 ;
        RECT 105.185 157.710 105.485 159.670 ;
        RECT 90.300 156.715 90.620 156.975 ;
        RECT 38.860 156.420 43.650 156.590 ;
        RECT 45.570 156.420 52.065 156.590 ;
        RECT 52.280 156.420 58.775 156.590 ;
        RECT 58.990 156.420 84.090 156.590 ;
        RECT 37.055 154.055 37.225 154.325 ;
        RECT 37.000 154.020 37.280 154.055 ;
        RECT 36.990 153.705 37.290 154.020 ;
        RECT 36.980 153.445 37.300 153.705 ;
        RECT 34.610 152.230 34.980 152.510 ;
        RECT 33.110 150.730 33.480 151.010 ;
        RECT 33.145 148.010 33.445 150.730 ;
        RECT 34.645 149.510 34.945 152.230 ;
        RECT 36.095 152.220 36.485 152.520 ;
        RECT 38.860 152.235 39.030 156.420 ;
        RECT 42.270 155.605 42.590 155.865 ;
        RECT 39.205 155.220 39.525 155.480 ;
        RECT 38.815 151.915 39.075 152.235 ;
        RECT 38.785 151.490 39.105 151.750 ;
        RECT 38.860 150.705 39.030 151.490 ;
        RECT 38.785 150.445 39.105 150.705 ;
        RECT 34.610 149.230 34.980 149.510 ;
        RECT 33.110 147.730 33.480 148.010 ;
        RECT 33.145 145.010 33.445 147.730 ;
        RECT 34.645 146.510 34.945 149.230 ;
        RECT 36.095 149.220 36.485 149.520 ;
        RECT 38.785 148.490 39.105 148.750 ;
        RECT 38.860 147.250 39.030 148.490 ;
        RECT 38.785 146.990 39.105 147.250 ;
        RECT 34.610 146.230 34.980 146.510 ;
        RECT 33.110 144.730 33.480 145.010 ;
        RECT 33.145 142.010 33.445 144.730 ;
        RECT 34.645 143.510 34.945 146.230 ;
        RECT 36.095 146.220 36.485 146.520 ;
        RECT 38.860 145.770 39.030 146.990 ;
        RECT 38.750 145.470 39.140 145.770 ;
        RECT 38.785 144.205 39.105 144.250 ;
        RECT 39.280 144.205 39.450 155.220 ;
        RECT 41.755 153.720 42.145 154.020 ;
        RECT 40.905 152.970 41.295 153.270 ;
        RECT 40.065 151.470 40.455 151.770 ;
        RECT 39.755 149.205 39.925 150.205 ;
        RECT 39.680 148.945 40.000 149.205 ;
        RECT 39.690 148.425 39.990 148.945 ;
        RECT 39.755 144.705 39.925 148.425 ;
        RECT 39.680 144.445 40.000 144.705 ;
        RECT 38.785 144.035 39.450 144.205 ;
        RECT 38.785 143.990 39.105 144.035 ;
        RECT 34.610 143.230 34.980 143.510 ;
        RECT 33.110 141.730 33.480 142.010 ;
        RECT 33.145 138.620 33.445 141.730 ;
        RECT 32.765 137.670 33.805 138.620 ;
        RECT 34.645 136.620 34.945 143.230 ;
        RECT 36.095 143.220 36.485 143.520 ;
        RECT 38.860 142.750 39.030 143.990 ;
        RECT 40.175 143.205 40.345 151.470 ;
        RECT 40.485 149.970 40.875 150.270 ;
        RECT 40.595 147.705 40.765 149.970 ;
        RECT 40.520 147.445 40.840 147.705 ;
        RECT 41.015 146.205 41.185 152.970 ;
        RECT 41.755 150.720 42.145 151.020 ;
        RECT 41.755 147.720 42.145 148.020 ;
        RECT 40.940 145.945 41.260 146.205 ;
        RECT 40.100 142.945 40.420 143.205 ;
        RECT 38.785 142.490 39.105 142.750 ;
        RECT 38.860 141.270 39.030 142.490 ;
        RECT 41.015 141.705 41.185 145.945 ;
        RECT 42.345 145.770 42.515 155.605 ;
        RECT 42.805 152.220 43.195 152.520 ;
        RECT 45.570 152.235 45.740 156.420 ;
        RECT 52.280 156.250 52.450 156.420 ;
        RECT 52.205 155.990 52.525 156.250 ;
        RECT 50.400 155.605 50.720 155.865 ;
        RECT 48.980 154.835 49.300 155.095 ;
        RECT 45.915 154.450 46.235 154.710 ;
        RECT 45.525 151.915 45.785 152.235 ;
        RECT 45.495 151.490 45.815 151.750 ;
        RECT 45.570 150.705 45.740 151.490 ;
        RECT 45.495 150.445 45.815 150.705 ;
        RECT 43.690 149.990 44.010 150.250 ;
        RECT 42.805 149.220 43.195 149.520 ;
        RECT 43.765 148.770 43.935 149.990 ;
        RECT 43.655 148.470 44.045 148.770 ;
        RECT 45.495 148.490 45.815 148.750 ;
        RECT 45.570 147.250 45.740 148.490 ;
        RECT 45.495 146.990 45.815 147.250 ;
        RECT 42.805 146.220 43.195 146.520 ;
        RECT 45.570 145.770 45.740 146.990 ;
        RECT 42.235 145.470 42.625 145.770 ;
        RECT 45.460 145.470 45.850 145.770 ;
        RECT 41.755 144.720 42.145 145.020 ;
        RECT 45.495 144.205 45.815 144.250 ;
        RECT 45.990 144.205 46.160 154.450 ;
        RECT 48.465 153.720 48.855 154.020 ;
        RECT 47.615 152.970 48.005 153.270 ;
        RECT 46.465 151.345 46.635 151.705 ;
        RECT 46.775 151.470 47.165 151.770 ;
        RECT 46.385 151.085 46.705 151.345 ;
        RECT 46.465 149.205 46.635 151.085 ;
        RECT 46.390 148.945 46.710 149.205 ;
        RECT 46.465 144.705 46.635 148.945 ;
        RECT 46.390 144.445 46.710 144.705 ;
        RECT 45.495 144.035 46.160 144.205 ;
        RECT 45.495 143.990 45.815 144.035 ;
        RECT 42.805 143.220 43.195 143.520 ;
        RECT 45.570 142.750 45.740 143.990 ;
        RECT 46.885 143.205 47.055 151.470 ;
        RECT 47.195 149.970 47.585 150.270 ;
        RECT 47.305 147.705 47.475 149.970 ;
        RECT 47.230 147.445 47.550 147.705 ;
        RECT 47.725 146.205 47.895 152.970 ;
        RECT 48.465 150.720 48.855 151.020 ;
        RECT 48.465 147.720 48.855 148.020 ;
        RECT 47.650 145.945 47.970 146.205 ;
        RECT 46.810 142.945 47.130 143.205 ;
        RECT 45.495 142.490 45.815 142.750 ;
        RECT 41.755 141.720 42.145 142.020 ;
        RECT 40.940 141.445 41.260 141.705 ;
        RECT 45.570 141.270 45.740 142.490 ;
        RECT 47.725 141.705 47.895 145.945 ;
        RECT 49.055 145.770 49.225 154.835 ;
        RECT 50.475 153.705 50.645 155.605 ;
        RECT 50.400 153.445 50.720 153.705 ;
        RECT 49.515 152.220 49.905 152.520 ;
        RECT 52.280 152.235 52.450 155.990 ;
        RECT 58.990 155.865 59.160 156.420 ;
        RECT 65.625 155.990 65.945 156.250 ;
        RECT 79.045 155.990 79.365 156.250 ;
        RECT 92.465 155.990 92.785 156.250 ;
        RECT 58.915 155.605 59.235 155.865 ;
        RECT 55.175 153.720 55.565 154.020 ;
        RECT 54.325 152.970 54.715 153.270 ;
        RECT 52.235 151.915 52.495 152.235 ;
        RECT 52.205 151.490 52.525 151.750 ;
        RECT 52.280 150.705 52.450 151.490 ;
        RECT 53.485 151.470 53.875 151.770 ;
        RECT 52.205 150.445 52.525 150.705 ;
        RECT 49.515 149.220 49.905 149.520 ;
        RECT 53.175 149.205 53.345 150.205 ;
        RECT 53.100 148.945 53.420 149.205 ;
        RECT 52.205 148.490 52.525 148.750 ;
        RECT 52.280 147.250 52.450 148.490 ;
        RECT 53.110 148.425 53.410 148.945 ;
        RECT 52.205 146.990 52.525 147.250 ;
        RECT 49.515 146.220 49.905 146.520 ;
        RECT 52.280 145.770 52.450 146.990 ;
        RECT 48.945 145.470 49.335 145.770 ;
        RECT 52.170 145.470 52.560 145.770 ;
        RECT 48.465 144.720 48.855 145.020 ;
        RECT 53.175 144.705 53.345 148.425 ;
        RECT 53.100 144.445 53.420 144.705 ;
        RECT 52.205 143.990 52.525 144.250 ;
        RECT 49.515 143.220 49.905 143.520 ;
        RECT 52.280 142.750 52.450 143.990 ;
        RECT 53.595 143.205 53.765 151.470 ;
        RECT 53.905 149.970 54.295 150.270 ;
        RECT 54.015 147.705 54.185 149.970 ;
        RECT 53.940 147.445 54.260 147.705 ;
        RECT 54.435 146.205 54.605 152.970 ;
        RECT 56.225 152.220 56.615 152.520 ;
        RECT 58.990 152.235 59.160 155.605 ;
        RECT 63.820 155.220 64.140 155.480 ;
        RECT 61.885 153.720 62.275 154.020 ;
        RECT 63.895 153.705 64.065 155.220 ;
        RECT 63.820 153.445 64.140 153.705 ;
        RECT 61.035 152.970 61.425 153.270 ;
        RECT 58.945 151.915 59.205 152.235 ;
        RECT 58.915 151.490 59.235 151.750 ;
        RECT 55.175 150.720 55.565 151.020 ;
        RECT 58.990 150.705 59.160 151.490 ;
        RECT 59.885 151.345 60.055 151.705 ;
        RECT 60.195 151.470 60.585 151.770 ;
        RECT 59.805 151.085 60.125 151.345 ;
        RECT 58.915 150.445 59.235 150.705 ;
        RECT 57.110 149.990 57.430 150.250 ;
        RECT 56.225 149.220 56.615 149.520 ;
        RECT 57.185 148.770 57.355 149.990 ;
        RECT 59.885 149.205 60.055 151.085 ;
        RECT 59.810 148.945 60.130 149.205 ;
        RECT 57.075 148.470 57.465 148.770 ;
        RECT 58.915 148.490 59.235 148.750 ;
        RECT 55.175 147.720 55.565 148.020 ;
        RECT 58.990 147.250 59.160 148.490 ;
        RECT 58.915 146.990 59.235 147.250 ;
        RECT 56.225 146.220 56.615 146.520 ;
        RECT 54.360 145.945 54.680 146.205 ;
        RECT 53.520 142.945 53.840 143.205 ;
        RECT 52.205 142.490 52.525 142.750 ;
        RECT 48.465 141.720 48.855 142.020 ;
        RECT 47.650 141.445 47.970 141.705 ;
        RECT 52.280 141.270 52.450 142.490 ;
        RECT 54.435 141.705 54.605 145.945 ;
        RECT 58.990 145.770 59.160 146.990 ;
        RECT 55.655 145.470 56.045 145.770 ;
        RECT 58.880 145.470 59.270 145.770 ;
        RECT 55.175 144.720 55.565 145.020 ;
        RECT 55.175 141.720 55.565 142.020 ;
        RECT 54.360 141.445 54.680 141.705 ;
        RECT 38.750 140.970 39.140 141.270 ;
        RECT 45.460 140.970 45.850 141.270 ;
        RECT 52.170 140.970 52.560 141.270 ;
        RECT 34.275 135.670 35.315 136.620 ;
        RECT 52.280 135.425 52.450 140.970 ;
        RECT 54.170 135.670 55.210 136.620 ;
        RECT 52.205 135.165 52.525 135.425 ;
        RECT 54.440 134.165 54.940 135.670 ;
        RECT 55.765 135.040 55.935 145.470 ;
        RECT 59.885 144.705 60.055 148.945 ;
        RECT 59.810 144.445 60.130 144.705 ;
        RECT 58.915 143.990 59.235 144.250 ;
        RECT 56.225 143.220 56.615 143.520 ;
        RECT 58.990 142.750 59.160 143.990 ;
        RECT 60.305 143.205 60.475 151.470 ;
        RECT 60.615 149.970 61.005 150.270 ;
        RECT 60.725 147.705 60.895 149.970 ;
        RECT 60.650 147.445 60.970 147.705 ;
        RECT 61.145 146.205 61.315 152.970 ;
        RECT 62.935 152.220 63.325 152.520 ;
        RECT 65.700 152.235 65.870 155.990 ;
        RECT 72.365 155.575 72.625 155.895 ;
        RECT 68.595 153.720 68.985 154.020 ;
        RECT 67.745 152.970 68.135 153.270 ;
        RECT 65.655 151.915 65.915 152.235 ;
        RECT 65.625 151.490 65.945 151.750 ;
        RECT 61.885 150.720 62.275 151.020 ;
        RECT 65.700 150.705 65.870 151.490 ;
        RECT 66.905 151.470 67.295 151.770 ;
        RECT 65.625 150.445 65.945 150.705 ;
        RECT 62.935 149.220 63.325 149.520 ;
        RECT 66.595 149.205 66.765 150.205 ;
        RECT 66.520 148.945 66.840 149.205 ;
        RECT 65.625 148.490 65.945 148.750 ;
        RECT 61.885 147.720 62.275 148.020 ;
        RECT 65.700 147.250 65.870 148.490 ;
        RECT 66.530 148.425 66.830 148.945 ;
        RECT 65.625 146.990 65.945 147.250 ;
        RECT 62.935 146.220 63.325 146.520 ;
        RECT 61.070 145.945 61.390 146.205 ;
        RECT 60.230 142.945 60.550 143.205 ;
        RECT 58.915 142.490 59.235 142.750 ;
        RECT 58.990 141.270 59.160 142.490 ;
        RECT 61.145 141.705 61.315 145.945 ;
        RECT 65.700 145.770 65.870 146.990 ;
        RECT 62.365 145.470 62.755 145.770 ;
        RECT 65.590 145.470 65.980 145.770 ;
        RECT 61.885 144.720 62.275 145.020 ;
        RECT 61.885 141.720 62.275 142.020 ;
        RECT 61.070 141.445 61.390 141.705 ;
        RECT 58.880 140.970 59.270 141.270 ;
        RECT 56.690 137.670 57.730 138.620 ;
        RECT 55.690 134.780 56.010 135.040 ;
        RECT 56.960 134.165 57.460 137.670 ;
        RECT 58.990 135.425 59.160 140.970 ;
        RECT 59.790 139.785 60.110 140.045 ;
        RECT 58.915 135.165 59.235 135.425 ;
        RECT 54.440 133.665 55.300 134.165 ;
        RECT 54.800 96.675 55.300 133.665 ;
        RECT 54.525 96.175 55.300 96.675 ;
        RECT 55.550 133.665 57.460 134.165 ;
        RECT 35.110 94.790 35.430 95.050 ;
        RECT 30.305 92.760 31.345 93.710 ;
        RECT 30.650 91.280 30.950 92.760 ;
        RECT 30.640 89.440 30.960 91.280 ;
        RECT 35.185 90.925 35.355 94.790 ;
        RECT 39.610 94.405 39.930 94.665 ;
        RECT 35.110 90.665 35.430 90.925 ;
        RECT 36.345 90.760 37.385 91.710 ;
        RECT 39.685 90.925 39.855 94.405 ;
        RECT 44.110 94.020 44.430 94.280 ;
        RECT 44.185 90.925 44.355 94.020 ;
        RECT 48.610 93.635 48.930 93.895 ;
        RECT 48.685 90.925 48.855 93.635 ;
        RECT 53.110 93.250 53.430 93.510 ;
        RECT 53.185 90.925 53.355 93.250 ;
        RECT 54.525 91.710 55.025 96.175 ;
        RECT 55.550 93.710 56.050 133.665 ;
        RECT 59.865 133.595 60.035 139.785 ;
        RECT 61.170 139.400 61.490 139.660 ;
        RECT 62.475 139.615 62.645 145.470 ;
        RECT 66.595 144.705 66.765 148.425 ;
        RECT 66.520 144.445 66.840 144.705 ;
        RECT 65.625 143.990 65.945 144.250 ;
        RECT 62.935 143.220 63.325 143.520 ;
        RECT 65.700 142.750 65.870 143.990 ;
        RECT 67.015 143.205 67.185 151.470 ;
        RECT 67.325 149.970 67.715 150.270 ;
        RECT 67.435 147.705 67.605 149.970 ;
        RECT 67.360 147.445 67.680 147.705 ;
        RECT 67.855 146.205 68.025 152.970 ;
        RECT 69.645 152.220 70.035 152.520 ;
        RECT 72.410 152.235 72.580 155.575 ;
        RECT 77.240 154.835 77.560 155.095 ;
        RECT 75.305 153.720 75.695 154.020 ;
        RECT 77.315 153.705 77.485 154.835 ;
        RECT 77.240 153.445 77.560 153.705 ;
        RECT 74.455 152.970 74.845 153.270 ;
        RECT 72.365 151.915 72.625 152.235 ;
        RECT 72.335 151.490 72.655 151.750 ;
        RECT 68.595 150.720 68.985 151.020 ;
        RECT 72.410 150.705 72.580 151.490 ;
        RECT 73.305 151.345 73.475 151.705 ;
        RECT 73.615 151.470 74.005 151.770 ;
        RECT 73.225 151.085 73.545 151.345 ;
        RECT 72.335 150.445 72.655 150.705 ;
        RECT 70.530 149.990 70.850 150.250 ;
        RECT 69.645 149.220 70.035 149.520 ;
        RECT 70.605 148.770 70.775 149.990 ;
        RECT 73.305 149.205 73.475 151.085 ;
        RECT 73.230 148.945 73.550 149.205 ;
        RECT 70.495 148.470 70.885 148.770 ;
        RECT 72.335 148.490 72.655 148.750 ;
        RECT 68.595 147.720 68.985 148.020 ;
        RECT 72.410 147.250 72.580 148.490 ;
        RECT 72.335 146.990 72.655 147.250 ;
        RECT 69.645 146.220 70.035 146.520 ;
        RECT 67.780 145.945 68.100 146.205 ;
        RECT 66.940 142.945 67.260 143.205 ;
        RECT 65.625 142.490 65.945 142.750 ;
        RECT 65.700 141.270 65.870 142.490 ;
        RECT 67.855 141.705 68.025 145.945 ;
        RECT 72.410 145.770 72.580 146.990 ;
        RECT 69.075 145.470 69.465 145.770 ;
        RECT 72.300 145.470 72.690 145.770 ;
        RECT 68.595 144.720 68.985 145.020 ;
        RECT 68.595 141.720 68.985 142.020 ;
        RECT 67.780 141.445 68.100 141.705 ;
        RECT 65.590 140.970 65.980 141.270 ;
        RECT 62.105 139.445 62.645 139.615 ;
        RECT 61.245 133.595 61.415 139.400 ;
        RECT 62.105 135.040 62.275 139.445 ;
        RECT 62.550 139.015 62.870 139.275 ;
        RECT 62.030 134.780 62.350 135.040 ;
        RECT 62.625 133.595 62.795 139.015 ;
        RECT 63.930 138.630 64.250 138.890 ;
        RECT 65.700 138.845 65.870 140.970 ;
        RECT 65.700 138.675 66.240 138.845 ;
        RECT 64.005 133.595 64.175 138.630 ;
        RECT 65.310 138.245 65.630 138.505 ;
        RECT 65.385 133.595 65.555 138.245 ;
        RECT 66.070 136.195 66.240 138.675 ;
        RECT 66.690 137.860 67.010 138.120 ;
        RECT 65.995 135.935 66.315 136.195 ;
        RECT 66.765 133.595 66.935 137.860 ;
        RECT 68.070 137.475 68.390 137.735 ;
        RECT 69.185 137.690 69.355 145.470 ;
        RECT 73.305 144.705 73.475 148.945 ;
        RECT 73.230 144.445 73.550 144.705 ;
        RECT 72.335 143.990 72.655 144.250 ;
        RECT 69.645 143.220 70.035 143.520 ;
        RECT 72.410 142.750 72.580 143.990 ;
        RECT 73.725 143.205 73.895 151.470 ;
        RECT 74.035 149.970 74.425 150.270 ;
        RECT 74.145 147.705 74.315 149.970 ;
        RECT 74.070 147.445 74.390 147.705 ;
        RECT 74.565 146.205 74.735 152.970 ;
        RECT 76.355 152.220 76.745 152.520 ;
        RECT 79.120 152.235 79.290 155.990 ;
        RECT 85.755 155.605 86.075 155.865 ;
        RECT 82.015 153.720 82.405 154.020 ;
        RECT 81.165 152.970 81.555 153.270 ;
        RECT 79.075 151.915 79.335 152.235 ;
        RECT 79.045 151.490 79.365 151.750 ;
        RECT 75.305 150.720 75.695 151.020 ;
        RECT 79.120 150.705 79.290 151.490 ;
        RECT 80.325 151.470 80.715 151.770 ;
        RECT 79.045 150.445 79.365 150.705 ;
        RECT 76.355 149.220 76.745 149.520 ;
        RECT 80.015 149.205 80.185 150.205 ;
        RECT 79.940 148.945 80.260 149.205 ;
        RECT 79.045 148.490 79.365 148.750 ;
        RECT 75.305 147.720 75.695 148.020 ;
        RECT 79.120 147.250 79.290 148.490 ;
        RECT 79.950 148.425 80.250 148.945 ;
        RECT 79.045 146.990 79.365 147.250 ;
        RECT 76.355 146.220 76.745 146.520 ;
        RECT 74.490 145.945 74.810 146.205 ;
        RECT 73.650 142.945 73.970 143.205 ;
        RECT 72.335 142.490 72.655 142.750 ;
        RECT 72.410 141.270 72.580 142.490 ;
        RECT 74.565 141.705 74.735 145.945 ;
        RECT 79.120 145.770 79.290 146.990 ;
        RECT 75.785 145.470 76.175 145.770 ;
        RECT 79.010 145.470 79.400 145.770 ;
        RECT 75.305 144.720 75.695 145.020 ;
        RECT 75.305 141.720 75.695 142.020 ;
        RECT 74.490 141.445 74.810 141.705 ;
        RECT 72.300 140.970 72.690 141.270 ;
        RECT 68.815 137.520 69.355 137.690 ;
        RECT 68.145 133.595 68.315 137.475 ;
        RECT 68.815 135.810 68.985 137.520 ;
        RECT 69.450 137.090 69.770 137.350 ;
        RECT 72.410 137.305 72.580 140.970 ;
        RECT 72.410 137.135 72.950 137.305 ;
        RECT 68.740 135.550 69.060 135.810 ;
        RECT 69.525 133.595 69.695 137.090 ;
        RECT 72.780 136.965 72.950 137.135 ;
        RECT 70.830 136.705 71.150 136.965 ;
        RECT 72.705 136.705 73.025 136.965 ;
        RECT 70.905 133.595 71.075 136.705 ;
        RECT 75.895 136.580 76.065 145.470 ;
        RECT 80.015 144.705 80.185 148.425 ;
        RECT 79.940 144.445 80.260 144.705 ;
        RECT 79.045 143.990 79.365 144.250 ;
        RECT 76.355 143.220 76.745 143.520 ;
        RECT 79.120 142.750 79.290 143.990 ;
        RECT 80.435 143.205 80.605 151.470 ;
        RECT 80.745 149.970 81.135 150.270 ;
        RECT 80.855 147.705 81.025 149.970 ;
        RECT 80.780 147.445 81.100 147.705 ;
        RECT 81.275 146.205 81.445 152.970 ;
        RECT 83.065 152.220 83.455 152.520 ;
        RECT 85.830 152.235 86.000 155.605 ;
        RECT 90.660 154.450 90.980 154.710 ;
        RECT 88.725 153.720 89.115 154.020 ;
        RECT 90.735 153.705 90.905 154.450 ;
        RECT 90.660 153.445 90.980 153.705 ;
        RECT 87.875 152.970 88.265 153.270 ;
        RECT 85.785 151.915 86.045 152.235 ;
        RECT 85.755 151.490 86.075 151.750 ;
        RECT 82.015 150.720 82.405 151.020 ;
        RECT 85.830 150.705 86.000 151.490 ;
        RECT 86.725 151.345 86.895 151.705 ;
        RECT 87.035 151.470 87.425 151.770 ;
        RECT 86.645 151.085 86.965 151.345 ;
        RECT 85.755 150.445 86.075 150.705 ;
        RECT 83.950 149.990 84.270 150.250 ;
        RECT 83.065 149.220 83.455 149.520 ;
        RECT 84.025 148.770 84.195 149.990 ;
        RECT 86.725 149.205 86.895 151.085 ;
        RECT 86.650 148.945 86.970 149.205 ;
        RECT 83.915 148.470 84.305 148.770 ;
        RECT 85.755 148.490 86.075 148.750 ;
        RECT 82.015 147.720 82.405 148.020 ;
        RECT 85.830 147.250 86.000 148.490 ;
        RECT 85.755 146.990 86.075 147.250 ;
        RECT 83.065 146.220 83.455 146.520 ;
        RECT 81.200 145.945 81.520 146.205 ;
        RECT 80.360 142.945 80.680 143.205 ;
        RECT 79.045 142.490 79.365 142.750 ;
        RECT 79.120 141.270 79.290 142.490 ;
        RECT 81.275 141.705 81.445 145.945 ;
        RECT 85.830 145.770 86.000 146.990 ;
        RECT 82.495 145.470 82.885 145.770 ;
        RECT 85.720 145.470 86.110 145.770 ;
        RECT 82.015 144.720 82.405 145.020 ;
        RECT 82.015 141.720 82.405 142.020 ;
        RECT 81.200 141.445 81.520 141.705 ;
        RECT 79.010 140.970 79.400 141.270 ;
        RECT 79.120 137.735 79.290 140.970 ;
        RECT 79.045 137.475 79.365 137.735 ;
        RECT 81.145 137.670 82.185 138.620 ;
        RECT 72.210 136.320 72.530 136.580 ;
        RECT 75.820 136.320 76.140 136.580 ;
        RECT 72.285 133.595 72.455 136.320 ;
        RECT 73.590 135.935 73.910 136.195 ;
        RECT 73.665 133.595 73.835 135.935 ;
        RECT 74.970 135.550 75.290 135.810 ;
        RECT 75.045 133.595 75.215 135.550 ;
        RECT 76.350 135.165 76.670 135.425 ;
        RECT 81.415 135.165 81.915 137.670 ;
        RECT 82.605 137.350 82.775 145.470 ;
        RECT 86.725 144.705 86.895 148.945 ;
        RECT 86.650 144.445 86.970 144.705 ;
        RECT 85.755 143.990 86.075 144.250 ;
        RECT 83.065 143.220 83.455 143.520 ;
        RECT 85.830 142.750 86.000 143.990 ;
        RECT 87.145 143.205 87.315 151.470 ;
        RECT 87.455 149.970 87.845 150.270 ;
        RECT 87.565 147.705 87.735 149.970 ;
        RECT 87.490 147.445 87.810 147.705 ;
        RECT 87.985 146.205 88.155 152.970 ;
        RECT 89.775 152.220 90.165 152.520 ;
        RECT 92.540 152.235 92.710 155.990 ;
        RECT 99.175 155.605 99.495 155.865 ;
        RECT 95.435 153.720 95.825 154.020 ;
        RECT 94.585 152.970 94.975 153.270 ;
        RECT 92.495 151.915 92.755 152.235 ;
        RECT 92.465 151.490 92.785 151.750 ;
        RECT 88.725 150.720 89.115 151.020 ;
        RECT 92.540 150.705 92.710 151.490 ;
        RECT 93.745 151.470 94.135 151.770 ;
        RECT 92.465 150.445 92.785 150.705 ;
        RECT 89.775 149.220 90.165 149.520 ;
        RECT 93.435 149.205 93.605 150.205 ;
        RECT 93.360 148.945 93.680 149.205 ;
        RECT 92.465 148.490 92.785 148.750 ;
        RECT 88.725 147.720 89.115 148.020 ;
        RECT 92.540 147.250 92.710 148.490 ;
        RECT 93.370 148.425 93.670 148.945 ;
        RECT 92.465 146.990 92.785 147.250 ;
        RECT 89.775 146.220 90.165 146.520 ;
        RECT 87.910 145.945 88.230 146.205 ;
        RECT 87.070 142.945 87.390 143.205 ;
        RECT 85.755 142.490 86.075 142.750 ;
        RECT 85.830 141.270 86.000 142.490 ;
        RECT 87.985 141.705 88.155 145.945 ;
        RECT 92.540 145.770 92.710 146.990 ;
        RECT 89.205 145.470 89.595 145.770 ;
        RECT 92.430 145.470 92.820 145.770 ;
        RECT 88.725 144.720 89.115 145.020 ;
        RECT 88.725 141.720 89.115 142.020 ;
        RECT 87.910 141.445 88.230 141.705 ;
        RECT 85.720 140.970 86.110 141.270 ;
        RECT 85.830 138.505 86.000 140.970 ;
        RECT 85.755 138.245 86.075 138.505 ;
        RECT 89.315 138.120 89.485 145.470 ;
        RECT 93.435 144.705 93.605 148.425 ;
        RECT 93.360 144.445 93.680 144.705 ;
        RECT 92.465 143.990 92.785 144.250 ;
        RECT 89.775 143.220 90.165 143.520 ;
        RECT 92.540 142.750 92.710 143.990 ;
        RECT 93.855 143.205 94.025 151.470 ;
        RECT 94.165 149.970 94.555 150.270 ;
        RECT 94.275 147.705 94.445 149.970 ;
        RECT 94.200 147.445 94.520 147.705 ;
        RECT 94.695 146.205 94.865 152.970 ;
        RECT 96.485 152.220 96.875 152.520 ;
        RECT 99.250 152.235 99.420 155.605 ;
        RECT 102.145 153.720 102.535 154.020 ;
        RECT 101.295 152.970 101.685 153.270 ;
        RECT 99.205 151.915 99.465 152.235 ;
        RECT 99.175 151.490 99.495 151.750 ;
        RECT 95.435 150.720 95.825 151.020 ;
        RECT 99.250 150.705 99.420 151.490 ;
        RECT 100.145 151.345 100.315 151.705 ;
        RECT 100.455 151.470 100.845 151.770 ;
        RECT 100.065 151.085 100.385 151.345 ;
        RECT 99.175 150.445 99.495 150.705 ;
        RECT 97.370 149.990 97.690 150.250 ;
        RECT 96.485 149.220 96.875 149.520 ;
        RECT 97.445 148.770 97.615 149.990 ;
        RECT 100.145 149.205 100.315 151.085 ;
        RECT 100.070 148.945 100.390 149.205 ;
        RECT 97.335 148.470 97.725 148.770 ;
        RECT 99.175 148.490 99.495 148.750 ;
        RECT 95.435 147.720 95.825 148.020 ;
        RECT 99.250 147.250 99.420 148.490 ;
        RECT 99.175 146.990 99.495 147.250 ;
        RECT 96.485 146.220 96.875 146.520 ;
        RECT 94.620 145.945 94.940 146.205 ;
        RECT 93.780 142.945 94.100 143.205 ;
        RECT 92.465 142.490 92.785 142.750 ;
        RECT 92.540 141.270 92.710 142.490 ;
        RECT 94.695 141.705 94.865 145.945 ;
        RECT 99.250 145.770 99.420 146.990 ;
        RECT 95.915 145.470 96.305 145.770 ;
        RECT 99.140 145.470 99.530 145.770 ;
        RECT 95.435 144.720 95.825 145.020 ;
        RECT 95.435 141.720 95.825 142.020 ;
        RECT 94.620 141.445 94.940 141.705 ;
        RECT 92.430 140.970 92.820 141.270 ;
        RECT 92.540 139.275 92.710 140.970 ;
        RECT 92.465 139.015 92.785 139.275 ;
        RECT 96.025 138.890 96.195 145.470 ;
        RECT 100.145 144.705 100.315 148.945 ;
        RECT 100.070 144.445 100.390 144.705 ;
        RECT 99.175 143.990 99.495 144.250 ;
        RECT 96.485 143.220 96.875 143.520 ;
        RECT 99.250 142.750 99.420 143.990 ;
        RECT 100.565 143.205 100.735 151.470 ;
        RECT 100.875 149.970 101.265 150.270 ;
        RECT 100.985 147.705 101.155 149.970 ;
        RECT 100.910 147.445 101.230 147.705 ;
        RECT 101.405 146.205 101.575 152.970 ;
        RECT 103.685 152.510 103.985 157.670 ;
        RECT 105.155 157.410 105.515 157.710 ;
        RECT 105.185 154.010 105.485 157.410 ;
        RECT 105.150 153.730 105.520 154.010 ;
        RECT 103.650 152.230 104.020 152.510 ;
        RECT 102.145 150.720 102.535 151.020 ;
        RECT 103.685 149.510 103.985 152.230 ;
        RECT 105.185 151.010 105.485 153.730 ;
        RECT 105.150 150.730 105.520 151.010 ;
        RECT 103.650 149.230 104.020 149.510 ;
        RECT 102.145 147.720 102.535 148.020 ;
        RECT 103.685 146.510 103.985 149.230 ;
        RECT 105.185 148.010 105.485 150.730 ;
        RECT 105.150 147.730 105.520 148.010 ;
        RECT 103.650 146.230 104.020 146.510 ;
        RECT 101.330 145.945 101.650 146.205 ;
        RECT 100.490 142.945 100.810 143.205 ;
        RECT 99.175 142.490 99.495 142.750 ;
        RECT 99.250 141.270 99.420 142.490 ;
        RECT 101.405 141.705 101.575 145.945 ;
        RECT 102.625 145.470 103.015 145.770 ;
        RECT 102.145 144.720 102.535 145.020 ;
        RECT 102.145 141.720 102.535 142.020 ;
        RECT 101.330 141.445 101.650 141.705 ;
        RECT 99.140 140.970 99.530 141.270 ;
        RECT 99.250 140.045 99.420 140.970 ;
        RECT 99.175 139.785 99.495 140.045 ;
        RECT 102.735 139.660 102.905 145.470 ;
        RECT 103.685 143.510 103.985 146.230 ;
        RECT 105.185 145.010 105.485 147.730 ;
        RECT 105.150 144.730 105.520 145.010 ;
        RECT 103.650 143.230 104.020 143.510 ;
        RECT 102.660 139.400 102.980 139.660 ;
        RECT 95.950 138.630 96.270 138.890 ;
        RECT 89.240 137.860 89.560 138.120 ;
        RECT 82.530 137.090 82.850 137.350 ;
        RECT 103.685 136.620 103.985 143.230 ;
        RECT 105.185 142.010 105.485 144.730 ;
        RECT 105.150 141.730 105.520 142.010 ;
        RECT 105.185 138.620 105.485 141.730 ;
        RECT 104.810 137.670 105.850 138.620 ;
        RECT 83.150 135.670 84.190 136.620 ;
        RECT 103.320 135.670 104.360 136.620 ;
        RECT 76.425 133.595 76.595 135.165 ;
        RECT 77.730 134.780 78.050 135.040 ;
        RECT 77.805 133.595 77.975 134.780 ;
        RECT 81.415 134.665 83.160 135.165 ;
        RECT 79.110 134.395 79.430 134.655 ;
        RECT 79.185 133.595 79.355 134.395 ;
        RECT 80.490 134.010 80.810 134.270 ;
        RECT 80.565 133.595 80.735 134.010 ;
        RECT 59.765 133.315 60.135 133.595 ;
        RECT 61.145 133.315 61.515 133.595 ;
        RECT 62.525 133.315 62.895 133.595 ;
        RECT 63.905 133.315 64.275 133.595 ;
        RECT 65.285 133.315 65.655 133.595 ;
        RECT 66.665 133.315 67.035 133.595 ;
        RECT 68.045 133.315 68.415 133.595 ;
        RECT 69.425 133.315 69.795 133.595 ;
        RECT 70.805 133.315 71.175 133.595 ;
        RECT 72.185 133.315 72.555 133.595 ;
        RECT 73.565 133.315 73.935 133.595 ;
        RECT 74.945 133.315 75.315 133.595 ;
        RECT 76.325 133.315 76.695 133.595 ;
        RECT 77.705 133.315 78.075 133.595 ;
        RECT 79.085 133.315 79.455 133.595 ;
        RECT 80.465 133.315 80.835 133.595 ;
        RECT 56.845 132.255 82.375 132.945 ;
        RECT 56.335 131.440 56.655 132.090 ;
        RECT 56.335 127.605 56.565 131.440 ;
        RECT 56.845 129.730 57.535 132.255 ;
        RECT 57.715 131.440 58.035 132.090 ;
        RECT 56.705 129.540 57.165 129.585 ;
        RECT 56.705 129.310 57.535 129.540 ;
        RECT 56.705 129.265 57.165 129.310 ;
        RECT 56.705 127.605 57.165 127.650 ;
        RECT 56.335 127.375 57.165 127.605 ;
        RECT 56.705 127.330 57.165 127.375 ;
        RECT 56.335 126.355 57.025 127.190 ;
        RECT 57.305 126.355 57.535 129.310 ;
        RECT 57.715 127.605 57.945 131.440 ;
        RECT 58.225 129.730 58.915 132.255 ;
        RECT 59.095 131.440 59.415 132.090 ;
        RECT 58.085 129.540 58.545 129.585 ;
        RECT 58.085 129.310 58.915 129.540 ;
        RECT 58.085 129.265 58.545 129.310 ;
        RECT 58.085 127.605 58.545 127.650 ;
        RECT 57.715 127.375 58.545 127.605 ;
        RECT 58.085 127.330 58.545 127.375 ;
        RECT 56.335 126.125 57.535 126.355 ;
        RECT 57.715 126.355 58.405 127.190 ;
        RECT 58.685 126.355 58.915 129.310 ;
        RECT 59.095 127.605 59.325 131.440 ;
        RECT 59.800 131.280 60.100 131.965 ;
        RECT 60.475 131.440 60.795 132.090 ;
        RECT 59.605 130.590 60.295 131.280 ;
        RECT 59.605 129.730 60.295 130.420 ;
        RECT 59.465 129.540 59.925 129.585 ;
        RECT 59.465 129.310 60.295 129.540 ;
        RECT 59.465 129.265 59.925 129.310 ;
        RECT 59.465 127.605 59.925 127.650 ;
        RECT 59.095 127.375 59.925 127.605 ;
        RECT 59.465 127.330 59.925 127.375 ;
        RECT 59.095 126.495 59.785 127.190 ;
        RECT 60.065 126.355 60.295 129.310 ;
        RECT 60.475 127.605 60.705 131.440 ;
        RECT 61.180 131.280 61.480 131.965 ;
        RECT 61.855 131.440 62.175 132.090 ;
        RECT 60.985 130.590 61.675 131.280 ;
        RECT 60.985 129.730 61.675 130.420 ;
        RECT 60.845 129.540 61.305 129.585 ;
        RECT 60.845 129.310 61.675 129.540 ;
        RECT 60.845 129.265 61.305 129.310 ;
        RECT 60.845 127.605 61.305 127.650 ;
        RECT 60.475 127.375 61.305 127.605 ;
        RECT 60.845 127.330 61.305 127.375 ;
        RECT 60.475 126.495 61.165 127.190 ;
        RECT 61.445 126.355 61.675 129.310 ;
        RECT 61.855 127.605 62.085 131.440 ;
        RECT 62.560 131.280 62.860 131.965 ;
        RECT 63.235 131.440 63.555 132.090 ;
        RECT 62.365 130.590 63.055 131.280 ;
        RECT 62.365 129.730 63.055 130.420 ;
        RECT 62.225 129.540 62.685 129.585 ;
        RECT 62.225 129.310 63.055 129.540 ;
        RECT 62.225 129.265 62.685 129.310 ;
        RECT 62.225 127.605 62.685 127.650 ;
        RECT 61.855 127.375 62.685 127.605 ;
        RECT 62.225 127.330 62.685 127.375 ;
        RECT 61.855 126.495 62.545 127.190 ;
        RECT 62.825 126.355 63.055 129.310 ;
        RECT 63.235 127.605 63.465 131.440 ;
        RECT 63.940 131.280 64.240 131.965 ;
        RECT 64.615 131.440 64.935 132.090 ;
        RECT 63.745 130.590 64.435 131.280 ;
        RECT 63.745 129.730 64.435 130.420 ;
        RECT 63.605 129.540 64.065 129.585 ;
        RECT 63.605 129.310 64.435 129.540 ;
        RECT 63.605 129.265 64.065 129.310 ;
        RECT 63.605 127.605 64.065 127.650 ;
        RECT 63.235 127.375 64.065 127.605 ;
        RECT 63.605 127.330 64.065 127.375 ;
        RECT 63.235 126.495 63.925 127.190 ;
        RECT 64.205 126.355 64.435 129.310 ;
        RECT 64.615 127.605 64.845 131.440 ;
        RECT 65.320 131.280 65.620 131.965 ;
        RECT 65.995 131.440 66.315 132.090 ;
        RECT 65.125 130.590 65.815 131.280 ;
        RECT 65.125 129.730 65.815 130.420 ;
        RECT 64.985 129.540 65.445 129.585 ;
        RECT 64.985 129.310 65.815 129.540 ;
        RECT 64.985 129.265 65.445 129.310 ;
        RECT 64.985 127.605 65.445 127.650 ;
        RECT 64.615 127.375 65.445 127.605 ;
        RECT 64.985 127.330 65.445 127.375 ;
        RECT 64.615 126.495 65.305 127.190 ;
        RECT 65.585 126.355 65.815 129.310 ;
        RECT 65.995 127.605 66.225 131.440 ;
        RECT 66.700 131.280 67.000 131.965 ;
        RECT 67.375 131.440 67.695 132.090 ;
        RECT 66.505 130.590 67.195 131.280 ;
        RECT 66.505 129.730 67.195 130.420 ;
        RECT 66.365 129.540 66.825 129.585 ;
        RECT 66.365 129.310 67.195 129.540 ;
        RECT 66.365 129.265 66.825 129.310 ;
        RECT 66.365 127.605 66.825 127.650 ;
        RECT 65.995 127.375 66.825 127.605 ;
        RECT 66.365 127.330 66.825 127.375 ;
        RECT 65.995 126.495 66.685 127.190 ;
        RECT 66.965 126.355 67.195 129.310 ;
        RECT 67.375 127.605 67.605 131.440 ;
        RECT 68.080 131.280 68.380 131.965 ;
        RECT 68.755 131.440 69.075 132.090 ;
        RECT 67.885 130.590 68.575 131.280 ;
        RECT 67.885 129.730 68.575 130.420 ;
        RECT 67.745 129.540 68.205 129.585 ;
        RECT 67.745 129.310 68.575 129.540 ;
        RECT 67.745 129.265 68.205 129.310 ;
        RECT 67.745 127.605 68.205 127.650 ;
        RECT 67.375 127.375 68.205 127.605 ;
        RECT 67.745 127.330 68.205 127.375 ;
        RECT 67.375 126.495 68.065 127.190 ;
        RECT 68.345 126.355 68.575 129.310 ;
        RECT 68.755 127.605 68.985 131.440 ;
        RECT 69.460 131.280 69.760 131.965 ;
        RECT 70.135 131.440 70.455 132.090 ;
        RECT 69.265 130.590 69.955 131.280 ;
        RECT 69.265 129.730 69.955 130.420 ;
        RECT 69.125 129.540 69.585 129.585 ;
        RECT 69.125 129.310 69.955 129.540 ;
        RECT 69.125 129.265 69.585 129.310 ;
        RECT 69.125 127.605 69.585 127.650 ;
        RECT 68.755 127.375 69.585 127.605 ;
        RECT 69.125 127.330 69.585 127.375 ;
        RECT 68.755 126.495 69.445 127.190 ;
        RECT 69.725 126.355 69.955 129.310 ;
        RECT 70.135 127.605 70.365 131.440 ;
        RECT 70.840 131.280 71.140 131.965 ;
        RECT 71.515 131.440 71.835 132.090 ;
        RECT 70.645 130.590 71.335 131.280 ;
        RECT 70.645 129.730 71.335 130.420 ;
        RECT 70.505 129.540 70.965 129.585 ;
        RECT 70.505 129.310 71.335 129.540 ;
        RECT 70.505 129.265 70.965 129.310 ;
        RECT 70.505 127.605 70.965 127.650 ;
        RECT 70.135 127.375 70.965 127.605 ;
        RECT 70.505 127.330 70.965 127.375 ;
        RECT 70.135 126.495 70.825 127.190 ;
        RECT 71.105 126.355 71.335 129.310 ;
        RECT 71.515 127.605 71.745 131.440 ;
        RECT 72.220 131.280 72.520 131.965 ;
        RECT 72.895 131.440 73.215 132.090 ;
        RECT 72.025 130.590 72.715 131.280 ;
        RECT 72.025 129.730 72.715 130.420 ;
        RECT 71.885 129.540 72.345 129.585 ;
        RECT 71.885 129.310 72.715 129.540 ;
        RECT 71.885 129.265 72.345 129.310 ;
        RECT 71.885 127.605 72.345 127.650 ;
        RECT 71.515 127.375 72.345 127.605 ;
        RECT 71.885 127.330 72.345 127.375 ;
        RECT 71.515 126.495 72.205 127.190 ;
        RECT 72.485 126.355 72.715 129.310 ;
        RECT 72.895 127.605 73.125 131.440 ;
        RECT 73.600 131.280 73.900 131.965 ;
        RECT 74.275 131.440 74.595 132.090 ;
        RECT 73.405 130.590 74.095 131.280 ;
        RECT 73.405 129.730 74.095 130.420 ;
        RECT 73.265 129.540 73.725 129.585 ;
        RECT 73.265 129.310 74.095 129.540 ;
        RECT 73.265 129.265 73.725 129.310 ;
        RECT 73.265 127.605 73.725 127.650 ;
        RECT 72.895 127.375 73.725 127.605 ;
        RECT 73.265 127.330 73.725 127.375 ;
        RECT 72.895 126.495 73.585 127.190 ;
        RECT 73.865 126.355 74.095 129.310 ;
        RECT 74.275 127.605 74.505 131.440 ;
        RECT 74.980 131.280 75.280 131.965 ;
        RECT 75.655 131.440 75.975 132.090 ;
        RECT 74.785 130.590 75.475 131.280 ;
        RECT 74.785 129.730 75.475 130.420 ;
        RECT 74.645 129.540 75.105 129.585 ;
        RECT 74.645 129.310 75.475 129.540 ;
        RECT 74.645 129.265 75.105 129.310 ;
        RECT 74.645 127.605 75.105 127.650 ;
        RECT 74.275 127.375 75.105 127.605 ;
        RECT 74.645 127.330 75.105 127.375 ;
        RECT 74.275 126.495 74.965 127.190 ;
        RECT 75.245 126.355 75.475 129.310 ;
        RECT 75.655 127.605 75.885 131.440 ;
        RECT 76.360 131.280 76.660 131.965 ;
        RECT 77.035 131.440 77.355 132.090 ;
        RECT 76.165 130.590 76.855 131.280 ;
        RECT 76.165 129.730 76.855 130.420 ;
        RECT 76.025 129.540 76.485 129.585 ;
        RECT 76.025 129.310 76.855 129.540 ;
        RECT 76.025 129.265 76.485 129.310 ;
        RECT 76.025 127.605 76.485 127.650 ;
        RECT 75.655 127.375 76.485 127.605 ;
        RECT 76.025 127.330 76.485 127.375 ;
        RECT 75.655 126.495 76.345 127.190 ;
        RECT 76.625 126.355 76.855 129.310 ;
        RECT 77.035 127.605 77.265 131.440 ;
        RECT 77.740 131.280 78.040 131.965 ;
        RECT 78.415 131.440 78.735 132.090 ;
        RECT 77.545 130.590 78.235 131.280 ;
        RECT 77.545 129.730 78.235 130.420 ;
        RECT 77.405 129.540 77.865 129.585 ;
        RECT 77.405 129.310 78.235 129.540 ;
        RECT 77.405 129.265 77.865 129.310 ;
        RECT 77.405 127.605 77.865 127.650 ;
        RECT 77.035 127.375 77.865 127.605 ;
        RECT 77.405 127.330 77.865 127.375 ;
        RECT 77.035 126.495 77.725 127.190 ;
        RECT 78.005 126.355 78.235 129.310 ;
        RECT 78.415 127.605 78.645 131.440 ;
        RECT 79.120 131.280 79.420 131.965 ;
        RECT 79.795 131.440 80.115 132.090 ;
        RECT 78.925 130.590 79.615 131.280 ;
        RECT 78.925 129.730 79.615 130.420 ;
        RECT 78.785 129.540 79.245 129.585 ;
        RECT 78.785 129.310 79.615 129.540 ;
        RECT 78.785 129.265 79.245 129.310 ;
        RECT 78.785 127.605 79.245 127.650 ;
        RECT 78.415 127.375 79.245 127.605 ;
        RECT 78.785 127.330 79.245 127.375 ;
        RECT 78.415 126.495 79.105 127.190 ;
        RECT 79.385 126.355 79.615 129.310 ;
        RECT 79.795 127.605 80.025 131.440 ;
        RECT 80.500 131.280 80.800 131.965 ;
        RECT 81.175 131.440 81.495 132.090 ;
        RECT 80.305 130.590 80.995 131.280 ;
        RECT 80.305 129.730 80.995 130.420 ;
        RECT 80.165 129.540 80.625 129.585 ;
        RECT 80.165 129.310 80.995 129.540 ;
        RECT 80.165 129.265 80.625 129.310 ;
        RECT 80.165 127.605 80.625 127.650 ;
        RECT 79.795 127.375 80.625 127.605 ;
        RECT 80.165 127.330 80.625 127.375 ;
        RECT 79.795 126.495 80.485 127.190 ;
        RECT 80.765 126.355 80.995 129.310 ;
        RECT 81.175 127.605 81.405 131.440 ;
        RECT 81.685 129.730 82.375 132.255 ;
        RECT 81.545 129.540 82.005 129.585 ;
        RECT 81.545 129.310 82.375 129.540 ;
        RECT 81.545 129.265 82.005 129.310 ;
        RECT 81.545 127.605 82.005 127.650 ;
        RECT 81.175 127.375 82.005 127.605 ;
        RECT 81.545 127.330 82.005 127.375 ;
        RECT 57.715 126.125 58.915 126.355 ;
        RECT 59.580 126.125 60.295 126.355 ;
        RECT 60.960 126.125 61.675 126.355 ;
        RECT 62.340 126.125 63.055 126.355 ;
        RECT 63.720 126.125 64.435 126.355 ;
        RECT 65.100 126.125 65.815 126.355 ;
        RECT 66.480 126.125 67.195 126.355 ;
        RECT 67.860 126.125 68.575 126.355 ;
        RECT 69.240 126.125 69.955 126.355 ;
        RECT 70.620 126.125 71.335 126.355 ;
        RECT 72.000 126.125 72.715 126.355 ;
        RECT 73.380 126.125 74.095 126.355 ;
        RECT 74.760 126.125 75.475 126.355 ;
        RECT 76.140 126.125 76.855 126.355 ;
        RECT 77.520 126.125 78.235 126.355 ;
        RECT 78.900 126.125 79.615 126.355 ;
        RECT 80.280 126.125 80.995 126.355 ;
        RECT 81.175 126.355 81.865 127.190 ;
        RECT 82.145 126.355 82.375 129.310 ;
        RECT 81.175 126.125 82.375 126.355 ;
        RECT 56.335 125.470 57.050 126.125 ;
        RECT 57.305 125.665 57.565 125.985 ;
        RECT 56.335 125.150 57.165 125.470 ;
        RECT 57.305 124.910 57.535 125.665 ;
        RECT 56.845 124.220 57.535 124.910 ;
        RECT 57.715 125.470 58.430 126.125 ;
        RECT 58.685 125.665 58.945 125.985 ;
        RECT 59.580 125.840 59.810 126.125 ;
        RECT 57.715 125.150 58.545 125.470 ;
        RECT 57.715 124.910 58.405 125.150 ;
        RECT 58.685 124.910 58.915 125.665 ;
        RECT 59.095 125.470 59.810 125.840 ;
        RECT 60.065 125.665 60.325 125.985 ;
        RECT 60.960 125.840 61.190 126.125 ;
        RECT 59.095 125.150 59.925 125.470 ;
        RECT 60.065 124.910 60.295 125.665 ;
        RECT 60.475 125.470 61.190 125.840 ;
        RECT 61.445 125.665 61.705 125.985 ;
        RECT 62.340 125.840 62.570 126.125 ;
        RECT 60.475 125.150 61.305 125.470 ;
        RECT 61.445 124.910 61.675 125.665 ;
        RECT 61.855 125.470 62.570 125.840 ;
        RECT 62.825 125.665 63.085 125.985 ;
        RECT 63.720 125.840 63.950 126.125 ;
        RECT 61.855 125.150 62.685 125.470 ;
        RECT 62.825 124.910 63.055 125.665 ;
        RECT 63.235 125.470 63.950 125.840 ;
        RECT 64.205 125.665 64.465 125.985 ;
        RECT 65.100 125.840 65.330 126.125 ;
        RECT 63.235 125.150 64.065 125.470 ;
        RECT 64.205 124.910 64.435 125.665 ;
        RECT 64.615 125.470 65.330 125.840 ;
        RECT 65.585 125.665 65.845 125.985 ;
        RECT 66.480 125.840 66.710 126.125 ;
        RECT 64.615 125.150 65.445 125.470 ;
        RECT 65.585 124.910 65.815 125.665 ;
        RECT 65.995 125.470 66.710 125.840 ;
        RECT 66.965 125.665 67.225 125.985 ;
        RECT 67.860 125.840 68.090 126.125 ;
        RECT 65.995 125.150 66.825 125.470 ;
        RECT 66.965 124.910 67.195 125.665 ;
        RECT 67.375 125.470 68.090 125.840 ;
        RECT 68.345 125.665 68.605 125.985 ;
        RECT 69.240 125.840 69.470 126.125 ;
        RECT 67.375 125.150 68.205 125.470 ;
        RECT 68.345 124.910 68.575 125.665 ;
        RECT 68.755 125.470 69.470 125.840 ;
        RECT 69.725 125.665 69.985 125.985 ;
        RECT 70.620 125.840 70.850 126.125 ;
        RECT 68.755 125.150 69.585 125.470 ;
        RECT 69.725 124.910 69.955 125.665 ;
        RECT 70.135 125.470 70.850 125.840 ;
        RECT 71.105 125.665 71.365 125.985 ;
        RECT 72.000 125.840 72.230 126.125 ;
        RECT 70.135 125.150 70.965 125.470 ;
        RECT 71.105 124.910 71.335 125.665 ;
        RECT 71.515 125.470 72.230 125.840 ;
        RECT 72.485 125.665 72.745 125.985 ;
        RECT 73.380 125.840 73.610 126.125 ;
        RECT 71.515 125.150 72.345 125.470 ;
        RECT 72.485 124.910 72.715 125.665 ;
        RECT 72.895 125.470 73.610 125.840 ;
        RECT 73.865 125.665 74.125 125.985 ;
        RECT 74.760 125.840 74.990 126.125 ;
        RECT 72.895 125.150 73.725 125.470 ;
        RECT 73.865 124.910 74.095 125.665 ;
        RECT 74.275 125.470 74.990 125.840 ;
        RECT 75.245 125.665 75.505 125.985 ;
        RECT 76.140 125.840 76.370 126.125 ;
        RECT 74.275 125.150 75.105 125.470 ;
        RECT 75.245 124.910 75.475 125.665 ;
        RECT 75.655 125.470 76.370 125.840 ;
        RECT 76.625 125.665 76.885 125.985 ;
        RECT 77.520 125.840 77.750 126.125 ;
        RECT 75.655 125.150 76.485 125.470 ;
        RECT 76.625 124.910 76.855 125.665 ;
        RECT 77.035 125.470 77.750 125.840 ;
        RECT 78.005 125.665 78.265 125.985 ;
        RECT 78.900 125.840 79.130 126.125 ;
        RECT 77.035 125.150 77.865 125.470 ;
        RECT 78.005 124.910 78.235 125.665 ;
        RECT 78.415 125.470 79.130 125.840 ;
        RECT 79.385 125.665 79.645 125.985 ;
        RECT 80.280 125.840 80.510 126.125 ;
        RECT 78.415 125.150 79.245 125.470 ;
        RECT 79.385 124.910 79.615 125.665 ;
        RECT 79.795 125.470 80.510 125.840 ;
        RECT 80.765 125.665 81.025 125.985 ;
        RECT 79.795 125.150 80.625 125.470 ;
        RECT 80.765 124.910 80.995 125.665 ;
        RECT 81.175 125.470 81.890 126.125 ;
        RECT 82.145 125.665 82.405 125.985 ;
        RECT 81.175 125.150 82.005 125.470 ;
        RECT 82.145 124.910 82.375 125.665 ;
        RECT 57.715 124.695 58.915 124.910 ;
        RECT 58.225 124.220 58.915 124.695 ;
        RECT 59.605 124.220 60.295 124.910 ;
        RECT 60.985 124.220 61.675 124.910 ;
        RECT 62.365 124.220 63.055 124.910 ;
        RECT 63.745 124.220 64.435 124.910 ;
        RECT 65.125 124.220 65.815 124.910 ;
        RECT 66.505 124.220 67.195 124.910 ;
        RECT 67.885 124.220 68.575 124.910 ;
        RECT 69.265 124.220 69.955 124.910 ;
        RECT 70.645 124.220 71.335 124.910 ;
        RECT 72.025 124.220 72.715 124.910 ;
        RECT 73.405 124.220 74.095 124.910 ;
        RECT 74.785 124.220 75.475 124.910 ;
        RECT 76.165 124.220 76.855 124.910 ;
        RECT 77.545 124.220 78.235 124.910 ;
        RECT 78.925 124.220 79.615 124.910 ;
        RECT 80.305 124.220 80.995 124.910 ;
        RECT 81.685 124.220 82.375 124.910 ;
        RECT 56.845 123.135 82.375 123.825 ;
        RECT 77.065 122.370 77.415 122.395 ;
        RECT 77.895 122.370 78.245 122.395 ;
        RECT 78.725 122.370 79.075 122.395 ;
        RECT 79.555 122.370 79.905 122.395 ;
        RECT 80.385 122.370 80.735 122.395 ;
        RECT 81.215 122.370 81.565 122.395 ;
        RECT 77.045 122.070 77.435 122.370 ;
        RECT 77.875 122.070 78.265 122.370 ;
        RECT 78.705 122.070 79.095 122.370 ;
        RECT 79.535 122.070 79.925 122.370 ;
        RECT 80.365 122.070 80.755 122.370 ;
        RECT 81.195 122.070 81.585 122.370 ;
        RECT 76.235 121.965 76.585 121.990 ;
        RECT 76.215 121.665 76.605 121.965 ;
        RECT 75.405 121.315 75.755 121.340 ;
        RECT 75.385 121.015 75.775 121.315 ;
        RECT 74.575 120.665 74.925 120.690 ;
        RECT 74.555 120.365 74.945 120.665 ;
        RECT 74.575 120.215 74.925 120.365 ;
        RECT 56.315 119.865 57.110 120.215 ;
        RECT 57.945 119.865 58.355 120.215 ;
        RECT 59.605 119.865 60.015 120.215 ;
        RECT 61.265 119.865 61.675 120.215 ;
        RECT 62.925 119.865 63.335 120.215 ;
        RECT 64.585 119.865 64.995 120.215 ;
        RECT 66.245 119.865 66.655 120.215 ;
        RECT 67.905 119.865 68.315 120.215 ;
        RECT 71.225 119.865 71.635 120.215 ;
        RECT 72.885 119.865 73.295 120.215 ;
        RECT 73.745 120.015 74.095 120.040 ;
        RECT 56.315 107.260 56.665 119.865 ;
        RECT 57.115 109.115 57.525 109.465 ;
        RECT 57.145 107.260 57.495 109.115 ;
        RECT 57.975 107.260 58.325 119.865 ;
        RECT 58.775 109.115 59.185 109.465 ;
        RECT 58.805 107.260 59.155 109.115 ;
        RECT 59.635 107.260 59.985 119.865 ;
        RECT 60.435 109.115 60.845 109.465 ;
        RECT 60.465 107.260 60.815 109.115 ;
        RECT 61.295 107.260 61.645 119.865 ;
        RECT 62.095 109.115 62.505 109.465 ;
        RECT 62.125 107.665 62.475 109.115 ;
        RECT 62.955 108.315 63.305 119.865 ;
        RECT 64.615 109.615 64.965 119.865 ;
        RECT 66.275 110.915 66.625 119.865 ;
        RECT 67.935 112.215 68.285 119.865 ;
        RECT 69.595 118.390 70.390 118.740 ;
        RECT 69.595 116.765 69.945 118.390 ;
        RECT 71.255 118.065 71.605 119.865 ;
        RECT 72.915 119.365 73.265 119.865 ;
        RECT 73.725 119.715 74.115 120.015 ;
        RECT 74.545 119.865 74.955 120.215 ;
        RECT 72.895 119.065 73.285 119.365 ;
        RECT 72.915 119.040 73.265 119.065 ;
        RECT 72.085 118.715 72.435 118.740 ;
        RECT 72.065 118.415 72.455 118.715 ;
        RECT 71.235 117.765 71.625 118.065 ;
        RECT 71.255 117.740 71.605 117.765 ;
        RECT 70.425 117.415 70.775 117.440 ;
        RECT 70.405 117.115 70.795 117.415 ;
        RECT 69.575 116.465 69.965 116.765 ;
        RECT 69.595 114.215 69.945 116.465 ;
        RECT 69.550 113.865 69.990 114.215 ;
        RECT 69.180 113.515 69.530 113.570 ;
        RECT 69.160 113.215 69.550 113.515 ;
        RECT 69.180 113.160 69.530 113.215 ;
        RECT 68.765 112.865 69.115 112.890 ;
        RECT 68.745 112.565 69.135 112.865 ;
        RECT 67.915 111.915 68.305 112.215 ;
        RECT 67.935 111.890 68.285 111.915 ;
        RECT 67.105 111.565 67.455 111.590 ;
        RECT 67.085 111.265 67.475 111.565 ;
        RECT 66.255 110.615 66.645 110.915 ;
        RECT 66.275 110.590 66.625 110.615 ;
        RECT 65.445 110.265 65.795 110.290 ;
        RECT 65.425 109.965 65.815 110.265 ;
        RECT 63.755 109.115 64.165 109.465 ;
        RECT 64.595 109.315 64.985 109.615 ;
        RECT 65.445 109.465 65.795 109.965 ;
        RECT 67.105 109.465 67.455 111.265 ;
        RECT 68.765 109.465 69.115 112.565 ;
        RECT 70.425 109.465 70.775 117.115 ;
        RECT 72.085 109.465 72.435 118.415 ;
        RECT 73.745 109.465 74.095 119.715 ;
        RECT 75.405 109.465 75.755 121.015 ;
        RECT 76.235 120.215 76.585 121.665 ;
        RECT 76.205 119.865 76.615 120.215 ;
        RECT 77.065 109.465 77.415 122.070 ;
        RECT 77.895 120.215 78.245 122.070 ;
        RECT 77.865 119.865 78.275 120.215 ;
        RECT 78.725 109.465 79.075 122.070 ;
        RECT 79.555 120.215 79.905 122.070 ;
        RECT 79.525 119.865 79.935 120.215 ;
        RECT 80.385 109.465 80.735 122.070 ;
        RECT 81.215 120.215 81.565 122.070 ;
        RECT 81.185 119.865 81.595 120.215 ;
        RECT 82.045 109.465 82.395 109.495 ;
        RECT 64.615 109.290 64.965 109.315 ;
        RECT 65.415 109.115 65.825 109.465 ;
        RECT 67.075 109.115 67.485 109.465 ;
        RECT 68.735 109.115 69.145 109.465 ;
        RECT 70.395 109.115 70.805 109.465 ;
        RECT 72.055 109.115 72.465 109.465 ;
        RECT 73.715 109.115 74.125 109.465 ;
        RECT 75.375 109.115 75.785 109.465 ;
        RECT 77.035 109.115 77.445 109.465 ;
        RECT 78.695 109.115 79.105 109.465 ;
        RECT 80.355 109.115 80.765 109.465 ;
        RECT 81.600 109.440 82.395 109.465 ;
        RECT 81.600 109.140 82.415 109.440 ;
        RECT 81.600 109.115 82.395 109.140 ;
        RECT 63.785 108.965 64.135 109.115 ;
        RECT 82.045 109.085 82.395 109.115 ;
        RECT 63.765 108.665 64.155 108.965 ;
        RECT 63.785 108.640 64.135 108.665 ;
        RECT 62.935 108.015 63.325 108.315 ;
        RECT 62.955 107.990 63.305 108.015 ;
        RECT 62.105 107.365 62.495 107.665 ;
        RECT 62.125 107.340 62.475 107.365 ;
        RECT 56.295 106.960 56.685 107.260 ;
        RECT 57.125 106.960 57.515 107.260 ;
        RECT 57.955 106.960 58.345 107.260 ;
        RECT 58.785 106.960 59.175 107.260 ;
        RECT 59.615 106.960 60.005 107.260 ;
        RECT 60.445 106.960 60.835 107.260 ;
        RECT 61.275 106.960 61.665 107.260 ;
        RECT 56.315 106.935 56.665 106.960 ;
        RECT 57.145 106.935 57.495 106.960 ;
        RECT 57.975 106.935 58.325 106.960 ;
        RECT 58.805 106.935 59.155 106.960 ;
        RECT 59.635 106.935 59.985 106.960 ;
        RECT 60.465 106.935 60.815 106.960 ;
        RECT 61.295 106.935 61.645 106.960 ;
        RECT 56.335 105.505 81.865 106.195 ;
        RECT 56.335 104.420 57.025 105.110 ;
        RECT 57.715 104.420 58.405 105.110 ;
        RECT 59.095 104.420 59.785 105.110 ;
        RECT 60.475 104.420 61.165 105.110 ;
        RECT 61.855 104.420 62.545 105.110 ;
        RECT 63.235 104.420 63.925 105.110 ;
        RECT 64.615 104.420 65.305 105.110 ;
        RECT 65.995 104.420 66.685 105.110 ;
        RECT 67.375 104.420 68.065 105.110 ;
        RECT 68.755 104.420 69.445 105.110 ;
        RECT 70.135 104.420 70.825 105.110 ;
        RECT 71.515 104.420 72.205 105.110 ;
        RECT 72.895 104.420 73.585 105.110 ;
        RECT 74.275 104.420 74.965 105.110 ;
        RECT 75.655 104.420 76.345 105.110 ;
        RECT 77.035 104.420 77.725 105.110 ;
        RECT 78.415 104.420 79.105 105.110 ;
        RECT 79.795 104.420 80.485 105.110 ;
        RECT 81.175 104.420 81.865 105.110 ;
        RECT 56.335 103.665 56.565 104.420 ;
        RECT 56.705 103.860 57.535 104.180 ;
        RECT 56.305 103.345 56.565 103.665 ;
        RECT 56.820 103.205 57.535 103.860 ;
        RECT 57.715 103.665 57.945 104.420 ;
        RECT 58.085 103.860 58.915 104.180 ;
        RECT 57.685 103.345 57.945 103.665 ;
        RECT 58.200 103.490 58.915 103.860 ;
        RECT 59.095 103.665 59.325 104.420 ;
        RECT 59.465 103.860 60.295 104.180 ;
        RECT 58.200 103.205 58.430 103.490 ;
        RECT 59.065 103.345 59.325 103.665 ;
        RECT 59.580 103.490 60.295 103.860 ;
        RECT 60.475 103.665 60.705 104.420 ;
        RECT 60.845 103.860 61.675 104.180 ;
        RECT 59.580 103.205 59.810 103.490 ;
        RECT 60.445 103.345 60.705 103.665 ;
        RECT 60.960 103.490 61.675 103.860 ;
        RECT 61.855 103.665 62.085 104.420 ;
        RECT 62.225 103.860 63.055 104.180 ;
        RECT 60.960 103.205 61.190 103.490 ;
        RECT 61.825 103.345 62.085 103.665 ;
        RECT 62.340 103.490 63.055 103.860 ;
        RECT 63.235 103.665 63.465 104.420 ;
        RECT 63.605 103.860 64.435 104.180 ;
        RECT 62.340 103.205 62.570 103.490 ;
        RECT 63.205 103.345 63.465 103.665 ;
        RECT 63.720 103.490 64.435 103.860 ;
        RECT 64.615 103.665 64.845 104.420 ;
        RECT 64.985 103.860 65.815 104.180 ;
        RECT 63.720 103.205 63.950 103.490 ;
        RECT 64.585 103.345 64.845 103.665 ;
        RECT 65.100 103.490 65.815 103.860 ;
        RECT 65.995 103.665 66.225 104.420 ;
        RECT 66.365 103.860 67.195 104.180 ;
        RECT 65.100 103.205 65.330 103.490 ;
        RECT 65.965 103.345 66.225 103.665 ;
        RECT 66.480 103.490 67.195 103.860 ;
        RECT 67.375 103.665 67.605 104.420 ;
        RECT 67.745 103.860 68.575 104.180 ;
        RECT 66.480 103.205 66.710 103.490 ;
        RECT 67.345 103.345 67.605 103.665 ;
        RECT 67.860 103.490 68.575 103.860 ;
        RECT 68.755 103.665 68.985 104.420 ;
        RECT 69.125 103.860 69.955 104.180 ;
        RECT 67.860 103.205 68.090 103.490 ;
        RECT 68.725 103.345 68.985 103.665 ;
        RECT 69.240 103.490 69.955 103.860 ;
        RECT 70.135 103.665 70.365 104.420 ;
        RECT 70.505 103.860 71.335 104.180 ;
        RECT 69.240 103.205 69.470 103.490 ;
        RECT 70.105 103.345 70.365 103.665 ;
        RECT 70.620 103.490 71.335 103.860 ;
        RECT 71.515 103.665 71.745 104.420 ;
        RECT 71.885 103.860 72.715 104.180 ;
        RECT 70.620 103.205 70.850 103.490 ;
        RECT 71.485 103.345 71.745 103.665 ;
        RECT 72.000 103.490 72.715 103.860 ;
        RECT 72.895 103.665 73.125 104.420 ;
        RECT 73.265 103.860 74.095 104.180 ;
        RECT 72.000 103.205 72.230 103.490 ;
        RECT 72.865 103.345 73.125 103.665 ;
        RECT 73.380 103.490 74.095 103.860 ;
        RECT 74.275 103.665 74.505 104.420 ;
        RECT 74.645 103.860 75.475 104.180 ;
        RECT 73.380 103.205 73.610 103.490 ;
        RECT 74.245 103.345 74.505 103.665 ;
        RECT 74.760 103.490 75.475 103.860 ;
        RECT 75.655 103.665 75.885 104.420 ;
        RECT 76.025 103.860 76.855 104.180 ;
        RECT 74.760 103.205 74.990 103.490 ;
        RECT 75.625 103.345 75.885 103.665 ;
        RECT 76.140 103.490 76.855 103.860 ;
        RECT 77.035 103.665 77.265 104.420 ;
        RECT 77.405 103.860 78.235 104.180 ;
        RECT 76.140 103.205 76.370 103.490 ;
        RECT 77.005 103.345 77.265 103.665 ;
        RECT 77.520 103.490 78.235 103.860 ;
        RECT 78.415 103.665 78.645 104.420 ;
        RECT 78.785 103.860 79.615 104.180 ;
        RECT 77.520 103.205 77.750 103.490 ;
        RECT 78.385 103.345 78.645 103.665 ;
        RECT 78.900 103.490 79.615 103.860 ;
        RECT 79.795 103.665 80.025 104.420 ;
        RECT 80.165 103.860 80.995 104.180 ;
        RECT 78.900 103.205 79.130 103.490 ;
        RECT 79.765 103.345 80.025 103.665 ;
        RECT 80.280 103.490 80.995 103.860 ;
        RECT 81.175 103.665 81.405 104.420 ;
        RECT 81.545 103.860 82.375 104.180 ;
        RECT 80.280 103.205 80.510 103.490 ;
        RECT 81.145 103.345 81.405 103.665 ;
        RECT 81.660 103.205 82.375 103.860 ;
        RECT 56.335 102.975 57.535 103.205 ;
        RECT 56.335 100.020 56.565 102.975 ;
        RECT 56.845 102.140 57.535 102.975 ;
        RECT 57.715 102.975 58.430 103.205 ;
        RECT 59.095 102.975 59.810 103.205 ;
        RECT 60.475 102.975 61.190 103.205 ;
        RECT 61.855 102.975 62.570 103.205 ;
        RECT 63.235 102.975 63.950 103.205 ;
        RECT 64.615 102.975 65.330 103.205 ;
        RECT 65.995 102.975 66.710 103.205 ;
        RECT 67.375 102.975 68.090 103.205 ;
        RECT 68.755 102.975 69.470 103.205 ;
        RECT 70.135 102.975 70.850 103.205 ;
        RECT 71.515 102.975 72.230 103.205 ;
        RECT 72.895 102.975 73.610 103.205 ;
        RECT 74.275 102.975 74.990 103.205 ;
        RECT 75.655 102.975 76.370 103.205 ;
        RECT 77.035 102.975 77.750 103.205 ;
        RECT 78.415 102.975 79.130 103.205 ;
        RECT 79.795 102.975 80.510 103.205 ;
        RECT 81.175 102.975 82.375 103.205 ;
        RECT 56.705 101.955 57.165 102.000 ;
        RECT 56.705 101.725 57.535 101.955 ;
        RECT 56.705 101.680 57.165 101.725 ;
        RECT 56.705 100.020 57.165 100.065 ;
        RECT 56.335 99.790 57.165 100.020 ;
        RECT 56.705 99.745 57.165 99.790 ;
        RECT 56.335 97.075 57.025 99.600 ;
        RECT 57.305 97.890 57.535 101.725 ;
        RECT 57.715 100.020 57.945 102.975 ;
        RECT 58.225 102.140 58.915 102.835 ;
        RECT 58.085 101.955 58.545 102.000 ;
        RECT 58.085 101.725 58.915 101.955 ;
        RECT 58.085 101.680 58.545 101.725 ;
        RECT 58.085 100.020 58.545 100.065 ;
        RECT 57.715 99.790 58.545 100.020 ;
        RECT 58.085 99.745 58.545 99.790 ;
        RECT 57.715 98.910 58.405 99.600 ;
        RECT 57.715 98.050 58.405 98.740 ;
        RECT 57.215 97.240 57.535 97.890 ;
        RECT 57.910 97.375 58.210 98.050 ;
        RECT 58.685 97.890 58.915 101.725 ;
        RECT 59.095 100.020 59.325 102.975 ;
        RECT 59.605 102.140 60.295 102.835 ;
        RECT 59.465 101.955 59.925 102.000 ;
        RECT 59.465 101.725 60.295 101.955 ;
        RECT 59.465 101.680 59.925 101.725 ;
        RECT 59.465 100.020 59.925 100.065 ;
        RECT 59.095 99.790 59.925 100.020 ;
        RECT 59.465 99.745 59.925 99.790 ;
        RECT 59.095 98.910 59.785 99.600 ;
        RECT 59.095 98.050 59.785 98.740 ;
        RECT 58.595 97.240 58.915 97.890 ;
        RECT 59.290 97.375 59.590 98.050 ;
        RECT 60.065 97.890 60.295 101.725 ;
        RECT 60.475 100.020 60.705 102.975 ;
        RECT 60.985 102.140 61.675 102.835 ;
        RECT 60.845 101.955 61.305 102.000 ;
        RECT 60.845 101.725 61.675 101.955 ;
        RECT 60.845 101.680 61.305 101.725 ;
        RECT 60.845 100.020 61.305 100.065 ;
        RECT 60.475 99.790 61.305 100.020 ;
        RECT 60.845 99.745 61.305 99.790 ;
        RECT 60.475 98.910 61.165 99.600 ;
        RECT 60.475 98.050 61.165 98.740 ;
        RECT 59.975 97.240 60.295 97.890 ;
        RECT 60.670 97.375 60.970 98.050 ;
        RECT 61.445 97.890 61.675 101.725 ;
        RECT 61.855 100.020 62.085 102.975 ;
        RECT 62.365 102.140 63.055 102.835 ;
        RECT 62.225 101.955 62.685 102.000 ;
        RECT 62.225 101.725 63.055 101.955 ;
        RECT 62.225 101.680 62.685 101.725 ;
        RECT 62.225 100.020 62.685 100.065 ;
        RECT 61.855 99.790 62.685 100.020 ;
        RECT 62.225 99.745 62.685 99.790 ;
        RECT 61.855 98.910 62.545 99.600 ;
        RECT 61.855 98.050 62.545 98.740 ;
        RECT 61.355 97.240 61.675 97.890 ;
        RECT 62.050 97.375 62.350 98.050 ;
        RECT 62.825 97.890 63.055 101.725 ;
        RECT 63.235 100.020 63.465 102.975 ;
        RECT 63.745 102.140 64.435 102.835 ;
        RECT 63.605 101.955 64.065 102.000 ;
        RECT 63.605 101.725 64.435 101.955 ;
        RECT 63.605 101.680 64.065 101.725 ;
        RECT 63.605 100.020 64.065 100.065 ;
        RECT 63.235 99.790 64.065 100.020 ;
        RECT 63.605 99.745 64.065 99.790 ;
        RECT 63.235 98.910 63.925 99.600 ;
        RECT 63.235 98.050 63.925 98.740 ;
        RECT 62.735 97.240 63.055 97.890 ;
        RECT 63.430 97.375 63.730 98.050 ;
        RECT 64.205 97.890 64.435 101.725 ;
        RECT 64.615 100.020 64.845 102.975 ;
        RECT 65.125 102.140 65.815 102.835 ;
        RECT 64.985 101.955 65.445 102.000 ;
        RECT 64.985 101.725 65.815 101.955 ;
        RECT 64.985 101.680 65.445 101.725 ;
        RECT 64.985 100.020 65.445 100.065 ;
        RECT 64.615 99.790 65.445 100.020 ;
        RECT 64.985 99.745 65.445 99.790 ;
        RECT 64.615 98.910 65.305 99.600 ;
        RECT 64.615 98.050 65.305 98.740 ;
        RECT 64.115 97.240 64.435 97.890 ;
        RECT 64.810 97.375 65.110 98.050 ;
        RECT 65.585 97.890 65.815 101.725 ;
        RECT 65.995 100.020 66.225 102.975 ;
        RECT 66.505 102.140 67.195 102.835 ;
        RECT 66.365 101.955 66.825 102.000 ;
        RECT 66.365 101.725 67.195 101.955 ;
        RECT 66.365 101.680 66.825 101.725 ;
        RECT 66.365 100.020 66.825 100.065 ;
        RECT 65.995 99.790 66.825 100.020 ;
        RECT 66.365 99.745 66.825 99.790 ;
        RECT 65.995 98.910 66.685 99.600 ;
        RECT 65.995 98.050 66.685 98.740 ;
        RECT 65.495 97.240 65.815 97.890 ;
        RECT 66.190 97.375 66.490 98.050 ;
        RECT 66.965 97.890 67.195 101.725 ;
        RECT 67.375 100.020 67.605 102.975 ;
        RECT 67.885 102.140 68.575 102.835 ;
        RECT 67.745 101.955 68.205 102.000 ;
        RECT 67.745 101.725 68.575 101.955 ;
        RECT 67.745 101.680 68.205 101.725 ;
        RECT 67.745 100.020 68.205 100.065 ;
        RECT 67.375 99.790 68.205 100.020 ;
        RECT 67.745 99.745 68.205 99.790 ;
        RECT 67.375 98.910 68.065 99.600 ;
        RECT 67.375 98.050 68.065 98.740 ;
        RECT 66.875 97.240 67.195 97.890 ;
        RECT 67.570 97.375 67.870 98.050 ;
        RECT 68.345 97.890 68.575 101.725 ;
        RECT 68.755 100.020 68.985 102.975 ;
        RECT 69.265 102.140 69.955 102.835 ;
        RECT 69.125 101.955 69.585 102.000 ;
        RECT 69.125 101.725 69.955 101.955 ;
        RECT 69.125 101.680 69.585 101.725 ;
        RECT 69.125 100.020 69.585 100.065 ;
        RECT 68.755 99.790 69.585 100.020 ;
        RECT 69.125 99.745 69.585 99.790 ;
        RECT 68.755 98.910 69.445 99.600 ;
        RECT 68.755 98.050 69.445 98.740 ;
        RECT 68.255 97.240 68.575 97.890 ;
        RECT 68.950 97.375 69.250 98.050 ;
        RECT 69.725 97.890 69.955 101.725 ;
        RECT 70.135 100.020 70.365 102.975 ;
        RECT 70.645 102.140 71.335 102.835 ;
        RECT 70.505 101.955 70.965 102.000 ;
        RECT 70.505 101.725 71.335 101.955 ;
        RECT 70.505 101.680 70.965 101.725 ;
        RECT 70.505 100.020 70.965 100.065 ;
        RECT 70.135 99.790 70.965 100.020 ;
        RECT 70.505 99.745 70.965 99.790 ;
        RECT 70.135 98.910 70.825 99.600 ;
        RECT 70.135 98.050 70.825 98.740 ;
        RECT 69.635 97.240 69.955 97.890 ;
        RECT 70.330 97.375 70.630 98.050 ;
        RECT 71.105 97.890 71.335 101.725 ;
        RECT 71.515 100.020 71.745 102.975 ;
        RECT 72.025 102.140 72.715 102.835 ;
        RECT 71.885 101.955 72.345 102.000 ;
        RECT 71.885 101.725 72.715 101.955 ;
        RECT 71.885 101.680 72.345 101.725 ;
        RECT 71.885 100.020 72.345 100.065 ;
        RECT 71.515 99.790 72.345 100.020 ;
        RECT 71.885 99.745 72.345 99.790 ;
        RECT 71.515 98.910 72.205 99.600 ;
        RECT 71.515 98.050 72.205 98.740 ;
        RECT 71.015 97.240 71.335 97.890 ;
        RECT 71.710 97.375 72.010 98.050 ;
        RECT 72.485 97.890 72.715 101.725 ;
        RECT 72.895 100.020 73.125 102.975 ;
        RECT 73.405 102.140 74.095 102.835 ;
        RECT 73.265 101.955 73.725 102.000 ;
        RECT 73.265 101.725 74.095 101.955 ;
        RECT 73.265 101.680 73.725 101.725 ;
        RECT 73.265 100.020 73.725 100.065 ;
        RECT 72.895 99.790 73.725 100.020 ;
        RECT 73.265 99.745 73.725 99.790 ;
        RECT 72.895 98.910 73.585 99.600 ;
        RECT 72.895 98.050 73.585 98.740 ;
        RECT 72.395 97.240 72.715 97.890 ;
        RECT 73.090 97.375 73.390 98.050 ;
        RECT 73.865 97.890 74.095 101.725 ;
        RECT 74.275 100.020 74.505 102.975 ;
        RECT 74.785 102.140 75.475 102.835 ;
        RECT 74.645 101.955 75.105 102.000 ;
        RECT 74.645 101.725 75.475 101.955 ;
        RECT 74.645 101.680 75.105 101.725 ;
        RECT 74.645 100.020 75.105 100.065 ;
        RECT 74.275 99.790 75.105 100.020 ;
        RECT 74.645 99.745 75.105 99.790 ;
        RECT 74.275 98.910 74.965 99.600 ;
        RECT 74.275 98.050 74.965 98.740 ;
        RECT 73.775 97.240 74.095 97.890 ;
        RECT 74.470 97.375 74.770 98.050 ;
        RECT 75.245 97.890 75.475 101.725 ;
        RECT 75.655 100.020 75.885 102.975 ;
        RECT 76.165 102.140 76.855 102.835 ;
        RECT 76.025 101.955 76.485 102.000 ;
        RECT 76.025 101.725 76.855 101.955 ;
        RECT 76.025 101.680 76.485 101.725 ;
        RECT 76.025 100.020 76.485 100.065 ;
        RECT 75.655 99.790 76.485 100.020 ;
        RECT 76.025 99.745 76.485 99.790 ;
        RECT 75.655 98.910 76.345 99.600 ;
        RECT 75.655 98.050 76.345 98.740 ;
        RECT 75.155 97.240 75.475 97.890 ;
        RECT 75.850 97.375 76.150 98.050 ;
        RECT 76.625 97.890 76.855 101.725 ;
        RECT 77.035 100.020 77.265 102.975 ;
        RECT 77.545 102.140 78.235 102.835 ;
        RECT 77.405 101.955 77.865 102.000 ;
        RECT 77.405 101.725 78.235 101.955 ;
        RECT 77.405 101.680 77.865 101.725 ;
        RECT 77.405 100.020 77.865 100.065 ;
        RECT 77.035 99.790 77.865 100.020 ;
        RECT 77.405 99.745 77.865 99.790 ;
        RECT 77.035 98.910 77.725 99.600 ;
        RECT 77.035 98.050 77.725 98.740 ;
        RECT 76.535 97.240 76.855 97.890 ;
        RECT 77.230 97.375 77.530 98.050 ;
        RECT 78.005 97.890 78.235 101.725 ;
        RECT 78.415 100.020 78.645 102.975 ;
        RECT 78.925 102.140 79.615 102.835 ;
        RECT 78.785 101.955 79.245 102.000 ;
        RECT 78.785 101.725 79.615 101.955 ;
        RECT 78.785 101.680 79.245 101.725 ;
        RECT 78.785 100.020 79.245 100.065 ;
        RECT 78.415 99.790 79.245 100.020 ;
        RECT 78.785 99.745 79.245 99.790 ;
        RECT 78.415 98.910 79.105 99.600 ;
        RECT 78.415 98.050 79.105 98.740 ;
        RECT 77.915 97.240 78.235 97.890 ;
        RECT 78.610 97.375 78.910 98.050 ;
        RECT 79.385 97.890 79.615 101.725 ;
        RECT 79.795 100.020 80.025 102.975 ;
        RECT 80.305 102.140 80.995 102.835 ;
        RECT 80.165 101.955 80.625 102.000 ;
        RECT 80.165 101.725 80.995 101.955 ;
        RECT 80.165 101.680 80.625 101.725 ;
        RECT 80.165 100.020 80.625 100.065 ;
        RECT 79.795 99.790 80.625 100.020 ;
        RECT 80.165 99.745 80.625 99.790 ;
        RECT 79.795 98.910 80.485 99.600 ;
        RECT 79.795 98.050 80.485 98.740 ;
        RECT 79.295 97.240 79.615 97.890 ;
        RECT 79.990 97.375 80.290 98.050 ;
        RECT 80.765 97.890 80.995 101.725 ;
        RECT 81.175 100.020 81.405 102.975 ;
        RECT 81.685 102.140 82.375 102.975 ;
        RECT 81.545 101.955 82.005 102.000 ;
        RECT 81.545 101.725 82.375 101.955 ;
        RECT 81.545 101.680 82.005 101.725 ;
        RECT 81.545 100.020 82.005 100.065 ;
        RECT 81.175 99.790 82.005 100.020 ;
        RECT 81.545 99.745 82.005 99.790 ;
        RECT 80.675 97.240 80.995 97.890 ;
        RECT 81.175 97.075 81.865 99.600 ;
        RECT 82.145 97.890 82.375 101.725 ;
        RECT 82.055 97.240 82.375 97.890 ;
        RECT 56.335 96.385 81.865 97.075 ;
        RECT 57.875 95.755 58.245 96.035 ;
        RECT 59.255 95.755 59.625 96.035 ;
        RECT 60.635 95.755 61.005 96.035 ;
        RECT 62.015 95.755 62.385 96.035 ;
        RECT 63.395 95.755 63.765 96.035 ;
        RECT 64.775 95.755 65.145 96.035 ;
        RECT 66.155 95.755 66.525 96.035 ;
        RECT 67.535 95.755 67.905 96.035 ;
        RECT 68.915 95.755 69.285 96.035 ;
        RECT 70.295 95.755 70.665 96.035 ;
        RECT 71.675 95.755 72.045 96.035 ;
        RECT 73.055 95.755 73.425 96.035 ;
        RECT 74.435 95.755 74.805 96.035 ;
        RECT 75.815 95.755 76.185 96.035 ;
        RECT 77.195 95.755 77.565 96.035 ;
        RECT 78.575 95.755 78.945 96.035 ;
        RECT 79.955 95.755 80.325 96.035 ;
        RECT 57.975 95.050 58.145 95.755 ;
        RECT 57.900 94.790 58.220 95.050 ;
        RECT 59.355 94.665 59.525 95.755 ;
        RECT 59.280 94.405 59.600 94.665 ;
        RECT 60.735 94.280 60.905 95.755 ;
        RECT 60.660 94.020 60.980 94.280 ;
        RECT 62.115 93.895 62.285 95.755 ;
        RECT 55.270 92.760 56.310 93.710 ;
        RECT 62.040 93.635 62.360 93.895 ;
        RECT 63.495 93.510 63.665 95.755 ;
        RECT 63.420 93.250 63.740 93.510 ;
        RECT 64.875 93.125 65.045 95.755 ;
        RECT 57.610 92.865 57.930 93.125 ;
        RECT 64.800 92.865 65.120 93.125 ;
        RECT 36.715 89.810 37.015 90.760 ;
        RECT 39.610 90.665 39.930 90.925 ;
        RECT 44.110 90.665 44.430 90.925 ;
        RECT 48.610 90.665 48.930 90.925 ;
        RECT 53.110 90.665 53.430 90.925 ;
        RECT 54.255 90.760 55.295 91.710 ;
        RECT 57.685 90.925 57.855 92.865 ;
        RECT 66.255 92.740 66.425 95.755 ;
        RECT 62.110 92.480 62.430 92.740 ;
        RECT 66.180 92.480 66.500 92.740 ;
        RECT 62.185 90.925 62.355 92.480 ;
        RECT 67.635 92.355 67.805 95.755 ;
        RECT 69.015 95.435 69.185 95.755 ;
        RECT 68.940 95.175 69.260 95.435 ;
        RECT 70.395 95.050 70.565 95.755 ;
        RECT 71.110 95.175 71.430 95.435 ;
        RECT 70.320 94.790 70.640 95.050 ;
        RECT 66.610 92.095 66.930 92.355 ;
        RECT 67.560 92.095 67.880 92.355 ;
        RECT 66.685 90.925 66.855 92.095 ;
        RECT 71.185 90.925 71.355 95.175 ;
        RECT 71.775 94.665 71.945 95.755 ;
        RECT 71.700 94.405 72.020 94.665 ;
        RECT 73.155 94.280 73.325 95.755 ;
        RECT 73.080 94.020 73.400 94.280 ;
        RECT 74.535 93.895 74.705 95.755 ;
        RECT 75.225 94.790 75.545 95.050 ;
        RECT 74.460 93.635 74.780 93.895 ;
        RECT 75.300 91.685 75.470 94.790 ;
        RECT 75.915 93.510 76.085 95.755 ;
        RECT 75.840 93.250 76.160 93.510 ;
        RECT 77.295 93.125 77.465 95.755 ;
        RECT 77.220 92.865 77.540 93.125 ;
        RECT 78.675 92.740 78.845 95.755 ;
        RECT 78.600 92.480 78.920 92.740 ;
        RECT 80.055 92.355 80.225 95.755 ;
        RECT 82.660 95.675 83.160 134.665 ;
        RECT 82.155 95.175 83.160 95.675 ;
        RECT 80.495 94.405 80.815 94.665 ;
        RECT 79.980 92.095 80.300 92.355 ;
        RECT 80.570 91.685 80.740 94.405 ;
        RECT 82.155 93.710 82.655 95.175 ;
        RECT 81.885 92.760 82.925 93.710 ;
        RECT 83.410 91.710 83.910 135.670 ;
        RECT 107.535 130.525 108.385 130.545 ;
        RECT 115.090 130.525 115.940 130.545 ;
        RECT 107.510 129.625 115.965 130.525 ;
        RECT 107.535 129.605 108.385 129.625 ;
        RECT 115.090 129.605 115.940 129.625 ;
        RECT 84.610 94.020 84.930 94.280 ;
        RECT 75.300 91.515 75.855 91.685 ;
        RECT 75.685 90.925 75.855 91.515 ;
        RECT 80.185 91.515 80.740 91.685 ;
        RECT 80.185 90.925 80.355 91.515 ;
        RECT 57.610 90.665 57.930 90.925 ;
        RECT 62.110 90.665 62.430 90.925 ;
        RECT 66.610 90.665 66.930 90.925 ;
        RECT 71.110 90.665 71.430 90.925 ;
        RECT 75.610 90.665 75.930 90.925 ;
        RECT 80.110 90.665 80.430 90.925 ;
        RECT 83.145 90.760 84.185 91.710 ;
        RECT 84.685 90.925 84.855 94.020 ;
        RECT 89.110 93.635 89.430 93.895 ;
        RECT 89.185 90.925 89.355 93.635 ;
        RECT 93.610 93.250 93.930 93.510 ;
        RECT 93.685 90.925 93.855 93.250 ;
        RECT 98.110 92.865 98.430 93.125 ;
        RECT 98.185 90.925 98.355 92.865 ;
        RECT 107.285 92.760 108.325 93.710 ;
        RECT 102.610 92.480 102.930 92.740 ;
        RECT 102.685 90.925 102.855 92.480 ;
        RECT 107.110 92.095 107.430 92.355 ;
        RECT 84.610 90.665 84.930 90.925 ;
        RECT 89.110 90.665 89.430 90.925 ;
        RECT 93.610 90.665 93.930 90.925 ;
        RECT 98.110 90.665 98.430 90.925 ;
        RECT 102.610 90.665 102.930 90.925 ;
        RECT 104.065 90.760 105.105 91.710 ;
        RECT 107.185 90.925 107.355 92.095 ;
        RECT 107.680 91.280 107.980 92.760 ;
        RECT 104.440 89.865 104.740 90.760 ;
        RECT 107.110 90.665 107.430 90.925 ;
        RECT 35.605 89.510 37.015 89.810 ;
        RECT 103.175 89.565 104.740 89.865 ;
        RECT 30.650 83.195 30.950 89.440 ;
        RECT 32.140 88.680 32.400 88.755 ;
        RECT 33.640 88.680 33.900 88.755 ;
        RECT 34.685 88.680 34.945 88.755 ;
        RECT 32.140 88.510 34.945 88.680 ;
        RECT 32.140 88.435 32.400 88.510 ;
        RECT 33.640 88.435 33.900 88.510 ;
        RECT 34.685 88.435 34.945 88.510 ;
        RECT 35.605 87.645 35.905 89.510 ;
        RECT 36.640 88.680 36.900 88.755 ;
        RECT 38.140 88.680 38.400 88.755 ;
        RECT 39.185 88.680 39.445 88.755 ;
        RECT 36.640 88.510 39.445 88.680 ;
        RECT 36.640 88.435 36.900 88.510 ;
        RECT 38.140 88.435 38.400 88.510 ;
        RECT 39.185 88.435 39.445 88.510 ;
        RECT 41.140 88.680 41.400 88.755 ;
        RECT 42.640 88.680 42.900 88.755 ;
        RECT 43.685 88.680 43.945 88.755 ;
        RECT 41.140 88.510 43.945 88.680 ;
        RECT 41.140 88.435 41.400 88.510 ;
        RECT 42.640 88.435 42.900 88.510 ;
        RECT 43.685 88.435 43.945 88.510 ;
        RECT 45.640 88.680 45.900 88.755 ;
        RECT 47.140 88.680 47.400 88.755 ;
        RECT 48.185 88.680 48.445 88.755 ;
        RECT 45.640 88.510 48.445 88.680 ;
        RECT 45.640 88.435 45.900 88.510 ;
        RECT 47.140 88.435 47.400 88.510 ;
        RECT 48.185 88.435 48.445 88.510 ;
        RECT 50.140 88.680 50.400 88.755 ;
        RECT 51.640 88.680 51.900 88.755 ;
        RECT 52.685 88.680 52.945 88.755 ;
        RECT 50.140 88.510 52.945 88.680 ;
        RECT 50.140 88.435 50.400 88.510 ;
        RECT 51.640 88.435 51.900 88.510 ;
        RECT 52.685 88.435 52.945 88.510 ;
        RECT 54.640 88.680 54.900 88.755 ;
        RECT 56.140 88.680 56.400 88.755 ;
        RECT 57.185 88.680 57.445 88.755 ;
        RECT 54.640 88.510 57.445 88.680 ;
        RECT 54.640 88.435 54.900 88.510 ;
        RECT 56.140 88.435 56.400 88.510 ;
        RECT 57.185 88.435 57.445 88.510 ;
        RECT 59.140 88.680 59.400 88.755 ;
        RECT 60.640 88.680 60.900 88.755 ;
        RECT 61.685 88.680 61.945 88.755 ;
        RECT 59.140 88.510 61.945 88.680 ;
        RECT 59.140 88.435 59.400 88.510 ;
        RECT 60.640 88.435 60.900 88.510 ;
        RECT 61.685 88.435 61.945 88.510 ;
        RECT 63.640 88.680 63.900 88.755 ;
        RECT 65.140 88.680 65.400 88.755 ;
        RECT 66.185 88.680 66.445 88.755 ;
        RECT 63.640 88.510 66.445 88.680 ;
        RECT 63.640 88.435 63.900 88.510 ;
        RECT 65.140 88.435 65.400 88.510 ;
        RECT 66.185 88.435 66.445 88.510 ;
        RECT 68.140 88.680 68.400 88.755 ;
        RECT 69.640 88.680 69.900 88.755 ;
        RECT 70.685 88.680 70.945 88.755 ;
        RECT 68.140 88.510 70.945 88.680 ;
        RECT 68.140 88.435 68.400 88.510 ;
        RECT 69.640 88.435 69.900 88.510 ;
        RECT 70.685 88.435 70.945 88.510 ;
        RECT 72.640 88.680 72.900 88.755 ;
        RECT 74.140 88.680 74.400 88.755 ;
        RECT 75.185 88.680 75.445 88.755 ;
        RECT 72.640 88.510 75.445 88.680 ;
        RECT 72.640 88.435 72.900 88.510 ;
        RECT 74.140 88.435 74.400 88.510 ;
        RECT 75.185 88.435 75.445 88.510 ;
        RECT 77.140 88.680 77.400 88.755 ;
        RECT 78.640 88.680 78.900 88.755 ;
        RECT 79.685 88.680 79.945 88.755 ;
        RECT 77.140 88.510 79.945 88.680 ;
        RECT 77.140 88.435 77.400 88.510 ;
        RECT 78.640 88.435 78.900 88.510 ;
        RECT 79.685 88.435 79.945 88.510 ;
        RECT 81.640 88.680 81.900 88.755 ;
        RECT 83.140 88.680 83.400 88.755 ;
        RECT 84.185 88.680 84.445 88.755 ;
        RECT 81.640 88.510 84.445 88.680 ;
        RECT 81.640 88.435 81.900 88.510 ;
        RECT 83.140 88.435 83.400 88.510 ;
        RECT 84.185 88.435 84.445 88.510 ;
        RECT 86.140 88.680 86.400 88.755 ;
        RECT 87.640 88.680 87.900 88.755 ;
        RECT 88.685 88.680 88.945 88.755 ;
        RECT 86.140 88.510 88.945 88.680 ;
        RECT 86.140 88.435 86.400 88.510 ;
        RECT 87.640 88.435 87.900 88.510 ;
        RECT 88.685 88.435 88.945 88.510 ;
        RECT 90.640 88.680 90.900 88.755 ;
        RECT 92.140 88.680 92.400 88.755 ;
        RECT 93.185 88.680 93.445 88.755 ;
        RECT 90.640 88.510 93.445 88.680 ;
        RECT 90.640 88.435 90.900 88.510 ;
        RECT 92.140 88.435 92.400 88.510 ;
        RECT 93.185 88.435 93.445 88.510 ;
        RECT 95.140 88.680 95.400 88.755 ;
        RECT 96.640 88.680 96.900 88.755 ;
        RECT 97.685 88.680 97.945 88.755 ;
        RECT 95.140 88.510 97.945 88.680 ;
        RECT 95.140 88.435 95.400 88.510 ;
        RECT 96.640 88.435 96.900 88.510 ;
        RECT 97.685 88.435 97.945 88.510 ;
        RECT 99.640 88.680 99.900 88.755 ;
        RECT 101.140 88.680 101.400 88.755 ;
        RECT 102.185 88.680 102.445 88.755 ;
        RECT 99.640 88.510 102.445 88.680 ;
        RECT 99.640 88.435 99.900 88.510 ;
        RECT 101.140 88.435 101.400 88.510 ;
        RECT 102.185 88.435 102.445 88.510 ;
        RECT 34.820 87.345 35.905 87.645 ;
        RECT 103.175 87.645 103.475 89.565 ;
        RECT 107.670 89.440 107.990 91.280 ;
        RECT 104.140 88.680 104.400 88.755 ;
        RECT 105.640 88.680 105.900 88.755 ;
        RECT 106.685 88.680 106.945 88.755 ;
        RECT 104.140 88.510 106.945 88.680 ;
        RECT 104.140 88.435 104.400 88.510 ;
        RECT 105.640 88.435 105.900 88.510 ;
        RECT 106.685 88.435 106.945 88.510 ;
        RECT 103.175 87.345 104.740 87.645 ;
        RECT 31.655 86.275 31.975 86.535 ;
        RECT 33.155 86.275 33.475 86.535 ;
        RECT 31.730 86.070 31.900 86.275 ;
        RECT 31.655 85.810 31.975 86.070 ;
        RECT 33.230 85.445 33.400 86.275 ;
        RECT 33.155 85.185 33.475 85.445 ;
        RECT 34.820 84.695 35.120 87.345 ;
        RECT 36.155 86.275 36.475 86.535 ;
        RECT 37.655 86.275 37.975 86.535 ;
        RECT 40.655 86.275 40.975 86.535 ;
        RECT 42.155 86.275 42.475 86.535 ;
        RECT 45.155 86.275 45.475 86.535 ;
        RECT 46.655 86.275 46.975 86.535 ;
        RECT 49.655 86.275 49.975 86.535 ;
        RECT 51.155 86.275 51.475 86.535 ;
        RECT 54.155 86.275 54.475 86.535 ;
        RECT 55.655 86.275 55.975 86.535 ;
        RECT 58.655 86.275 58.975 86.535 ;
        RECT 60.155 86.275 60.475 86.535 ;
        RECT 63.155 86.275 63.475 86.535 ;
        RECT 64.655 86.275 64.975 86.535 ;
        RECT 67.655 86.275 67.975 86.535 ;
        RECT 69.155 86.275 69.475 86.535 ;
        RECT 72.155 86.275 72.475 86.535 ;
        RECT 73.655 86.275 73.975 86.535 ;
        RECT 76.655 86.275 76.975 86.535 ;
        RECT 78.155 86.275 78.475 86.535 ;
        RECT 81.155 86.275 81.475 86.535 ;
        RECT 82.655 86.275 82.975 86.535 ;
        RECT 85.655 86.275 85.975 86.535 ;
        RECT 87.155 86.275 87.475 86.535 ;
        RECT 90.155 86.275 90.475 86.535 ;
        RECT 91.655 86.275 91.975 86.535 ;
        RECT 94.655 86.275 94.975 86.535 ;
        RECT 96.155 86.275 96.475 86.535 ;
        RECT 99.155 86.275 99.475 86.535 ;
        RECT 100.655 86.275 100.975 86.535 ;
        RECT 103.655 86.275 103.975 86.535 ;
        RECT 36.230 85.445 36.400 86.275 ;
        RECT 36.155 85.185 36.475 85.445 ;
        RECT 37.730 85.060 37.900 86.275 ;
        RECT 40.730 85.060 40.900 86.275 ;
        RECT 37.655 84.800 37.975 85.060 ;
        RECT 40.655 84.800 40.975 85.060 ;
        RECT 34.790 84.395 35.150 84.695 ;
        RECT 42.230 84.675 42.400 86.275 ;
        RECT 45.230 84.675 45.400 86.275 ;
        RECT 42.155 84.415 42.475 84.675 ;
        RECT 45.155 84.415 45.475 84.675 ;
        RECT 30.650 82.895 33.620 83.195 ;
        RECT 33.320 77.595 33.620 82.895 ;
        RECT 33.285 77.315 33.655 77.595 ;
        RECT 33.320 74.595 33.620 77.315 ;
        RECT 34.820 76.095 35.120 84.395 ;
        RECT 46.730 84.290 46.900 86.275 ;
        RECT 49.730 84.290 49.900 86.275 ;
        RECT 46.655 84.030 46.975 84.290 ;
        RECT 49.655 84.030 49.975 84.290 ;
        RECT 51.230 83.905 51.400 86.275 ;
        RECT 54.230 83.905 54.400 86.275 ;
        RECT 51.155 83.645 51.475 83.905 ;
        RECT 54.155 83.645 54.475 83.905 ;
        RECT 55.730 83.520 55.900 86.275 ;
        RECT 58.730 83.520 58.900 86.275 ;
        RECT 55.655 83.260 55.975 83.520 ;
        RECT 58.655 83.260 58.975 83.520 ;
        RECT 60.230 83.135 60.400 86.275 ;
        RECT 63.230 83.135 63.400 86.275 ;
        RECT 60.155 82.875 60.475 83.135 ;
        RECT 62.665 82.875 62.985 83.135 ;
        RECT 63.155 82.875 63.475 83.135 ;
        RECT 55.955 82.105 56.275 82.365 ;
        RECT 49.245 81.335 49.565 81.595 ;
        RECT 42.535 80.565 42.855 80.825 ;
        RECT 35.825 79.795 36.145 80.055 ;
        RECT 34.785 75.815 35.155 76.095 ;
        RECT 33.285 74.315 33.655 74.595 ;
        RECT 33.320 71.595 33.620 74.315 ;
        RECT 34.820 73.095 35.120 75.815 ;
        RECT 35.900 73.855 36.070 79.795 ;
        RECT 39.310 79.410 39.630 79.670 ;
        RECT 39.385 78.355 39.555 79.410 ;
        RECT 39.275 78.055 39.665 78.355 ;
        RECT 37.155 77.620 37.475 77.880 ;
        RECT 36.270 77.305 36.660 77.605 ;
        RECT 36.270 74.305 36.660 74.605 ;
        RECT 35.790 73.555 36.180 73.855 ;
        RECT 37.230 73.380 37.400 77.620 ;
        RECT 39.385 76.835 39.555 78.055 ;
        RECT 39.310 76.575 39.630 76.835 ;
        RECT 37.995 76.120 38.315 76.380 ;
        RECT 37.155 73.120 37.475 73.380 ;
        RECT 34.785 72.815 35.155 73.095 ;
        RECT 33.285 71.315 33.655 71.595 ;
        RECT 33.320 68.595 33.620 71.315 ;
        RECT 34.820 70.095 35.120 72.815 ;
        RECT 36.270 71.305 36.660 71.605 ;
        RECT 34.785 69.815 35.155 70.095 ;
        RECT 33.285 68.315 33.655 68.595 ;
        RECT 33.320 65.595 33.620 68.315 ;
        RECT 34.820 67.095 35.120 69.815 ;
        RECT 36.270 68.305 36.660 68.605 ;
        RECT 34.785 66.815 35.155 67.095 ;
        RECT 33.285 65.315 33.655 65.595 ;
        RECT 33.320 63.710 33.620 65.315 ;
        RECT 32.940 62.760 33.980 63.710 ;
        RECT 34.820 61.710 35.120 66.815 ;
        RECT 37.230 66.355 37.400 73.120 ;
        RECT 37.575 71.620 37.895 71.880 ;
        RECT 37.650 69.355 37.820 71.620 ;
        RECT 37.540 69.055 37.930 69.355 ;
        RECT 38.070 67.855 38.240 76.120 ;
        RECT 39.385 75.335 39.555 76.575 ;
        RECT 41.930 75.805 42.320 76.105 ;
        RECT 39.310 75.075 39.630 75.335 ;
        RECT 38.415 74.620 38.735 74.880 ;
        RECT 38.490 70.380 38.660 74.620 ;
        RECT 42.610 73.855 42.780 80.565 ;
        RECT 46.020 80.180 46.340 80.440 ;
        RECT 46.095 78.355 46.265 80.180 ;
        RECT 45.985 78.055 46.375 78.355 ;
        RECT 43.865 77.620 44.185 77.880 ;
        RECT 42.980 77.305 43.370 77.605 ;
        RECT 42.980 74.305 43.370 74.605 ;
        RECT 39.275 73.555 39.665 73.855 ;
        RECT 42.500 73.555 42.890 73.855 ;
        RECT 39.385 72.335 39.555 73.555 ;
        RECT 43.940 73.380 44.110 77.620 ;
        RECT 46.095 76.835 46.265 78.055 ;
        RECT 46.020 76.575 46.340 76.835 ;
        RECT 44.705 76.120 45.025 76.380 ;
        RECT 43.865 73.120 44.185 73.380 ;
        RECT 41.930 72.805 42.320 73.105 ;
        RECT 39.310 72.075 39.630 72.335 ;
        RECT 39.385 70.835 39.555 72.075 ;
        RECT 42.980 71.305 43.370 71.605 ;
        RECT 39.310 70.575 39.630 70.835 ;
        RECT 41.080 70.555 41.470 70.855 ;
        RECT 38.415 70.120 38.735 70.380 ;
        RECT 38.490 68.240 38.660 70.120 ;
        RECT 41.190 69.335 41.360 70.555 ;
        RECT 41.930 69.805 42.320 70.105 ;
        RECT 41.115 69.075 41.435 69.335 ;
        RECT 39.310 68.620 39.630 68.880 ;
        RECT 38.420 67.980 38.740 68.240 ;
        RECT 37.960 67.555 38.350 67.855 ;
        RECT 38.490 67.620 38.660 67.980 ;
        RECT 39.385 67.835 39.555 68.620 ;
        RECT 42.980 68.305 43.370 68.605 ;
        RECT 39.310 67.575 39.630 67.835 ;
        RECT 39.340 67.090 39.600 67.410 ;
        RECT 37.120 66.055 37.510 66.355 ;
        RECT 36.270 65.305 36.660 65.605 ;
        RECT 39.385 63.720 39.555 67.090 ;
        RECT 41.930 66.805 42.320 67.105 ;
        RECT 43.940 66.355 44.110 73.120 ;
        RECT 44.285 71.620 44.605 71.880 ;
        RECT 44.360 69.355 44.530 71.620 ;
        RECT 44.250 69.055 44.640 69.355 ;
        RECT 44.780 67.855 44.950 76.120 ;
        RECT 46.095 75.335 46.265 76.575 ;
        RECT 48.640 75.805 49.030 76.105 ;
        RECT 46.020 75.075 46.340 75.335 ;
        RECT 45.125 74.620 45.445 74.880 ;
        RECT 45.200 70.900 45.370 74.620 ;
        RECT 49.320 73.855 49.490 81.335 ;
        RECT 52.730 80.950 53.050 81.210 ;
        RECT 52.805 78.355 52.975 80.950 ;
        RECT 52.695 78.055 53.085 78.355 ;
        RECT 50.575 77.620 50.895 77.880 ;
        RECT 49.690 77.305 50.080 77.605 ;
        RECT 49.690 74.305 50.080 74.605 ;
        RECT 45.985 73.555 46.375 73.855 ;
        RECT 49.210 73.555 49.600 73.855 ;
        RECT 46.095 72.335 46.265 73.555 ;
        RECT 50.650 73.380 50.820 77.620 ;
        RECT 52.805 76.835 52.975 78.055 ;
        RECT 52.730 76.575 53.050 76.835 ;
        RECT 51.415 76.120 51.735 76.380 ;
        RECT 50.575 73.120 50.895 73.380 ;
        RECT 48.640 72.805 49.030 73.105 ;
        RECT 46.020 72.075 46.340 72.335 ;
        RECT 45.135 70.380 45.435 70.900 ;
        RECT 46.095 70.835 46.265 72.075 ;
        RECT 49.690 71.305 50.080 71.605 ;
        RECT 46.020 70.575 46.340 70.835 ;
        RECT 45.125 70.120 45.445 70.380 ;
        RECT 45.200 69.120 45.370 70.120 ;
        RECT 48.640 69.805 49.030 70.105 ;
        RECT 46.020 68.620 46.340 68.880 ;
        RECT 44.670 67.555 45.060 67.855 ;
        RECT 46.095 67.835 46.265 68.620 ;
        RECT 49.690 68.305 50.080 68.605 ;
        RECT 46.020 67.575 46.340 67.835 ;
        RECT 46.050 67.090 46.310 67.410 ;
        RECT 43.830 66.055 44.220 66.355 ;
        RECT 42.980 65.305 43.370 65.605 ;
        RECT 39.310 63.460 39.630 63.720 ;
        RECT 46.095 63.335 46.265 67.090 ;
        RECT 48.640 66.805 49.030 67.105 ;
        RECT 50.650 66.355 50.820 73.120 ;
        RECT 50.995 71.620 51.315 71.880 ;
        RECT 51.070 69.355 51.240 71.620 ;
        RECT 50.960 69.055 51.350 69.355 ;
        RECT 51.490 67.855 51.660 76.120 ;
        RECT 52.805 75.335 52.975 76.575 ;
        RECT 55.350 75.805 55.740 76.105 ;
        RECT 52.730 75.075 53.050 75.335 ;
        RECT 51.835 74.620 52.155 74.880 ;
        RECT 51.910 70.380 52.080 74.620 ;
        RECT 56.030 73.855 56.200 82.105 ;
        RECT 59.440 81.720 59.760 81.980 ;
        RECT 59.515 78.355 59.685 81.720 ;
        RECT 59.405 78.055 59.795 78.355 ;
        RECT 57.285 77.620 57.605 77.880 ;
        RECT 56.400 77.305 56.790 77.605 ;
        RECT 56.400 74.305 56.790 74.605 ;
        RECT 52.695 73.555 53.085 73.855 ;
        RECT 55.920 73.555 56.310 73.855 ;
        RECT 52.805 72.335 52.975 73.555 ;
        RECT 57.360 73.380 57.530 77.620 ;
        RECT 59.515 76.835 59.685 78.055 ;
        RECT 59.440 76.575 59.760 76.835 ;
        RECT 58.125 76.120 58.445 76.380 ;
        RECT 57.285 73.120 57.605 73.380 ;
        RECT 55.350 72.805 55.740 73.105 ;
        RECT 52.730 72.075 53.050 72.335 ;
        RECT 52.805 70.835 52.975 72.075 ;
        RECT 56.400 71.305 56.790 71.605 ;
        RECT 52.730 70.575 53.050 70.835 ;
        RECT 54.500 70.555 54.890 70.855 ;
        RECT 51.835 70.120 52.155 70.380 ;
        RECT 51.910 68.240 52.080 70.120 ;
        RECT 54.610 69.335 54.780 70.555 ;
        RECT 55.350 69.805 55.740 70.105 ;
        RECT 54.535 69.075 54.855 69.335 ;
        RECT 52.730 68.620 53.050 68.880 ;
        RECT 51.840 67.980 52.160 68.240 ;
        RECT 51.380 67.555 51.770 67.855 ;
        RECT 51.910 67.620 52.080 67.980 ;
        RECT 52.805 67.835 52.975 68.620 ;
        RECT 56.400 68.305 56.790 68.605 ;
        RECT 52.730 67.575 53.050 67.835 ;
        RECT 52.760 67.090 53.020 67.410 ;
        RECT 50.540 66.055 50.930 66.355 ;
        RECT 47.825 65.620 48.145 65.880 ;
        RECT 47.900 64.875 48.070 65.620 ;
        RECT 49.690 65.305 50.080 65.605 ;
        RECT 47.825 64.615 48.145 64.875 ;
        RECT 52.805 63.720 52.975 67.090 ;
        RECT 55.350 66.805 55.740 67.105 ;
        RECT 57.360 66.355 57.530 73.120 ;
        RECT 57.705 71.620 58.025 71.880 ;
        RECT 57.780 69.355 57.950 71.620 ;
        RECT 57.670 69.055 58.060 69.355 ;
        RECT 58.200 67.855 58.370 76.120 ;
        RECT 59.515 75.335 59.685 76.575 ;
        RECT 62.060 75.805 62.450 76.105 ;
        RECT 59.440 75.075 59.760 75.335 ;
        RECT 58.545 74.620 58.865 74.880 ;
        RECT 58.620 70.900 58.790 74.620 ;
        RECT 62.740 73.855 62.910 82.875 ;
        RECT 64.730 82.750 64.900 86.275 ;
        RECT 67.730 82.750 67.900 86.275 ;
        RECT 64.655 82.490 64.975 82.750 ;
        RECT 66.150 82.490 66.470 82.750 ;
        RECT 67.655 82.490 67.975 82.750 ;
        RECT 66.225 78.355 66.395 82.490 ;
        RECT 69.230 82.365 69.400 86.275 ;
        RECT 69.875 83.645 70.195 83.905 ;
        RECT 69.155 82.105 69.475 82.365 ;
        RECT 69.950 80.780 70.120 83.645 ;
        RECT 72.230 82.365 72.400 86.275 ;
        RECT 72.860 83.260 73.180 83.520 ;
        RECT 72.155 82.105 72.475 82.365 ;
        RECT 69.450 80.610 70.120 80.780 ;
        RECT 66.115 78.055 66.505 78.355 ;
        RECT 63.995 77.620 64.315 77.880 ;
        RECT 63.110 77.305 63.500 77.605 ;
        RECT 63.110 74.305 63.500 74.605 ;
        RECT 59.405 73.555 59.795 73.855 ;
        RECT 62.630 73.555 63.020 73.855 ;
        RECT 59.515 72.335 59.685 73.555 ;
        RECT 64.070 73.380 64.240 77.620 ;
        RECT 66.225 76.835 66.395 78.055 ;
        RECT 66.150 76.575 66.470 76.835 ;
        RECT 64.835 76.120 65.155 76.380 ;
        RECT 63.995 73.120 64.315 73.380 ;
        RECT 62.060 72.805 62.450 73.105 ;
        RECT 59.440 72.075 59.760 72.335 ;
        RECT 58.555 70.380 58.855 70.900 ;
        RECT 59.515 70.835 59.685 72.075 ;
        RECT 63.110 71.305 63.500 71.605 ;
        RECT 59.440 70.575 59.760 70.835 ;
        RECT 58.545 70.120 58.865 70.380 ;
        RECT 58.620 69.120 58.790 70.120 ;
        RECT 62.060 69.805 62.450 70.105 ;
        RECT 59.440 68.620 59.760 68.880 ;
        RECT 58.090 67.555 58.480 67.855 ;
        RECT 59.515 67.835 59.685 68.620 ;
        RECT 63.110 68.305 63.500 68.605 ;
        RECT 59.440 67.575 59.760 67.835 ;
        RECT 59.470 67.090 59.730 67.410 ;
        RECT 57.250 66.055 57.640 66.355 ;
        RECT 56.400 65.305 56.790 65.605 ;
        RECT 52.730 63.460 53.050 63.720 ;
        RECT 59.515 63.335 59.685 67.090 ;
        RECT 62.060 66.805 62.450 67.105 ;
        RECT 64.070 66.355 64.240 73.120 ;
        RECT 64.415 71.620 64.735 71.880 ;
        RECT 64.490 69.355 64.660 71.620 ;
        RECT 64.380 69.055 64.770 69.355 ;
        RECT 64.910 67.855 65.080 76.120 ;
        RECT 66.225 75.335 66.395 76.575 ;
        RECT 68.770 75.805 69.160 76.105 ;
        RECT 66.150 75.075 66.470 75.335 ;
        RECT 65.255 74.620 65.575 74.880 ;
        RECT 65.330 70.380 65.500 74.620 ;
        RECT 69.450 73.855 69.620 80.610 ;
        RECT 72.935 78.355 73.105 83.260 ;
        RECT 73.730 81.980 73.900 86.275 ;
        RECT 76.085 84.415 76.405 84.675 ;
        RECT 73.655 81.720 73.975 81.980 ;
        RECT 72.825 78.055 73.215 78.355 ;
        RECT 70.705 77.620 71.025 77.880 ;
        RECT 69.820 77.305 70.210 77.605 ;
        RECT 69.820 74.305 70.210 74.605 ;
        RECT 66.115 73.555 66.505 73.855 ;
        RECT 69.340 73.555 69.730 73.855 ;
        RECT 66.225 72.335 66.395 73.555 ;
        RECT 70.780 73.380 70.950 77.620 ;
        RECT 72.935 76.835 73.105 78.055 ;
        RECT 72.860 76.575 73.180 76.835 ;
        RECT 71.545 76.120 71.865 76.380 ;
        RECT 70.705 73.120 71.025 73.380 ;
        RECT 68.770 72.805 69.160 73.105 ;
        RECT 66.150 72.075 66.470 72.335 ;
        RECT 66.225 70.835 66.395 72.075 ;
        RECT 69.820 71.305 70.210 71.605 ;
        RECT 66.150 70.575 66.470 70.835 ;
        RECT 67.920 70.555 68.310 70.855 ;
        RECT 65.255 70.120 65.575 70.380 ;
        RECT 65.330 68.240 65.500 70.120 ;
        RECT 68.030 69.335 68.200 70.555 ;
        RECT 68.770 69.805 69.160 70.105 ;
        RECT 67.955 69.075 68.275 69.335 ;
        RECT 66.150 68.620 66.470 68.880 ;
        RECT 65.260 67.980 65.580 68.240 ;
        RECT 64.800 67.555 65.190 67.855 ;
        RECT 65.330 67.620 65.500 67.980 ;
        RECT 66.225 67.835 66.395 68.620 ;
        RECT 69.820 68.305 70.210 68.605 ;
        RECT 66.150 67.575 66.470 67.835 ;
        RECT 66.180 67.090 66.440 67.410 ;
        RECT 63.960 66.055 64.350 66.355 ;
        RECT 61.245 65.620 61.565 65.880 ;
        RECT 61.320 64.490 61.490 65.620 ;
        RECT 63.110 65.305 63.500 65.605 ;
        RECT 61.245 64.230 61.565 64.490 ;
        RECT 66.225 63.750 66.395 67.090 ;
        RECT 68.770 66.805 69.160 67.105 ;
        RECT 70.780 66.355 70.950 73.120 ;
        RECT 71.125 71.620 71.445 71.880 ;
        RECT 71.200 69.355 71.370 71.620 ;
        RECT 71.090 69.055 71.480 69.355 ;
        RECT 71.620 67.855 71.790 76.120 ;
        RECT 72.935 75.335 73.105 76.575 ;
        RECT 75.480 75.805 75.870 76.105 ;
        RECT 72.860 75.075 73.180 75.335 ;
        RECT 71.965 74.620 72.285 74.880 ;
        RECT 72.040 70.900 72.210 74.620 ;
        RECT 76.160 73.855 76.330 84.415 ;
        RECT 76.730 81.980 76.900 86.275 ;
        RECT 76.655 81.720 76.975 81.980 ;
        RECT 78.230 81.595 78.400 86.275 ;
        RECT 79.570 84.030 79.890 84.290 ;
        RECT 78.155 81.335 78.475 81.595 ;
        RECT 79.645 78.355 79.815 84.030 ;
        RECT 81.230 81.595 81.400 86.275 ;
        RECT 81.155 81.335 81.475 81.595 ;
        RECT 82.730 81.210 82.900 86.275 ;
        RECT 83.295 85.185 83.615 85.445 ;
        RECT 82.655 80.950 82.975 81.210 ;
        RECT 83.370 80.780 83.540 85.185 ;
        RECT 85.730 81.210 85.900 86.275 ;
        RECT 86.280 84.800 86.600 85.060 ;
        RECT 85.655 80.950 85.975 81.210 ;
        RECT 82.870 80.610 83.540 80.780 ;
        RECT 79.535 78.055 79.925 78.355 ;
        RECT 77.415 77.620 77.735 77.880 ;
        RECT 76.530 77.305 76.920 77.605 ;
        RECT 76.530 74.305 76.920 74.605 ;
        RECT 72.825 73.555 73.215 73.855 ;
        RECT 76.050 73.555 76.440 73.855 ;
        RECT 72.935 72.335 73.105 73.555 ;
        RECT 77.490 73.380 77.660 77.620 ;
        RECT 79.645 76.835 79.815 78.055 ;
        RECT 79.570 76.575 79.890 76.835 ;
        RECT 78.255 76.120 78.575 76.380 ;
        RECT 77.415 73.120 77.735 73.380 ;
        RECT 75.480 72.805 75.870 73.105 ;
        RECT 72.860 72.075 73.180 72.335 ;
        RECT 71.975 70.380 72.275 70.900 ;
        RECT 72.935 70.835 73.105 72.075 ;
        RECT 76.530 71.305 76.920 71.605 ;
        RECT 72.860 70.575 73.180 70.835 ;
        RECT 71.965 70.120 72.285 70.380 ;
        RECT 72.040 69.120 72.210 70.120 ;
        RECT 75.480 69.805 75.870 70.105 ;
        RECT 72.860 68.620 73.180 68.880 ;
        RECT 71.510 67.555 71.900 67.855 ;
        RECT 72.935 67.835 73.105 68.620 ;
        RECT 76.530 68.305 76.920 68.605 ;
        RECT 72.860 67.575 73.180 67.835 ;
        RECT 72.890 67.090 73.150 67.410 ;
        RECT 70.670 66.055 71.060 66.355 ;
        RECT 69.820 65.305 70.210 65.605 ;
        RECT 66.180 63.430 66.440 63.750 ;
        RECT 72.935 63.335 73.105 67.090 ;
        RECT 75.480 66.805 75.870 67.105 ;
        RECT 77.490 66.355 77.660 73.120 ;
        RECT 77.835 71.620 78.155 71.880 ;
        RECT 77.910 69.355 78.080 71.620 ;
        RECT 77.800 69.055 78.190 69.355 ;
        RECT 78.330 67.855 78.500 76.120 ;
        RECT 79.645 75.335 79.815 76.575 ;
        RECT 82.190 75.805 82.580 76.105 ;
        RECT 79.570 75.075 79.890 75.335 ;
        RECT 78.675 74.620 78.995 74.880 ;
        RECT 78.750 70.380 78.920 74.620 ;
        RECT 82.870 73.855 83.040 80.610 ;
        RECT 86.355 78.355 86.525 84.800 ;
        RECT 87.230 80.825 87.400 86.275 ;
        RECT 90.230 80.825 90.400 86.275 ;
        RECT 87.155 80.565 87.475 80.825 ;
        RECT 90.155 80.565 90.475 80.825 ;
        RECT 91.730 80.440 91.900 86.275 ;
        RECT 94.730 80.440 94.900 86.275 ;
        RECT 91.655 80.180 91.975 80.440 ;
        RECT 94.655 80.180 94.975 80.440 ;
        RECT 96.230 80.055 96.400 86.275 ;
        RECT 99.230 80.055 99.400 86.275 ;
        RECT 96.155 79.795 96.475 80.055 ;
        RECT 99.155 79.795 99.475 80.055 ;
        RECT 100.730 79.670 100.900 86.275 ;
        RECT 103.730 79.670 103.900 86.275 ;
        RECT 104.440 85.210 104.740 87.345 ;
        RECT 105.155 86.275 105.475 86.535 ;
        RECT 105.230 86.070 105.400 86.275 ;
        RECT 105.155 85.810 105.475 86.070 ;
        RECT 104.440 84.910 105.660 85.210 ;
        RECT 105.360 84.695 105.660 84.910 ;
        RECT 105.330 84.395 105.690 84.695 ;
        RECT 100.655 79.410 100.975 79.670 ;
        RECT 103.655 79.410 103.975 79.670 ;
        RECT 86.245 78.055 86.635 78.355 ;
        RECT 92.955 78.055 93.345 78.355 ;
        RECT 99.665 78.055 100.055 78.355 ;
        RECT 84.125 77.620 84.445 77.880 ;
        RECT 83.240 77.305 83.630 77.605 ;
        RECT 83.240 74.305 83.630 74.605 ;
        RECT 79.535 73.555 79.925 73.855 ;
        RECT 82.760 73.555 83.150 73.855 ;
        RECT 79.645 72.335 79.815 73.555 ;
        RECT 84.200 73.380 84.370 77.620 ;
        RECT 86.355 76.835 86.525 78.055 ;
        RECT 90.835 77.620 91.155 77.880 ;
        RECT 89.950 77.305 90.340 77.605 ;
        RECT 86.280 76.575 86.600 76.835 ;
        RECT 84.965 76.120 85.285 76.380 ;
        RECT 84.125 73.120 84.445 73.380 ;
        RECT 82.190 72.805 82.580 73.105 ;
        RECT 79.570 72.075 79.890 72.335 ;
        RECT 79.645 70.835 79.815 72.075 ;
        RECT 83.240 71.305 83.630 71.605 ;
        RECT 79.570 70.575 79.890 70.835 ;
        RECT 81.340 70.555 81.730 70.855 ;
        RECT 78.675 70.120 78.995 70.380 ;
        RECT 78.750 68.240 78.920 70.120 ;
        RECT 81.450 69.335 81.620 70.555 ;
        RECT 82.190 69.805 82.580 70.105 ;
        RECT 81.375 69.075 81.695 69.335 ;
        RECT 79.570 68.620 79.890 68.880 ;
        RECT 78.680 67.980 79.000 68.240 ;
        RECT 78.220 67.555 78.610 67.855 ;
        RECT 78.750 67.620 78.920 67.980 ;
        RECT 79.645 67.835 79.815 68.620 ;
        RECT 83.240 68.305 83.630 68.605 ;
        RECT 79.570 67.575 79.890 67.835 ;
        RECT 79.600 67.090 79.860 67.410 ;
        RECT 77.380 66.055 77.770 66.355 ;
        RECT 74.665 65.620 74.985 65.880 ;
        RECT 74.740 64.105 74.910 65.620 ;
        RECT 76.530 65.305 76.920 65.605 ;
        RECT 74.665 63.845 74.985 64.105 ;
        RECT 79.645 63.720 79.815 67.090 ;
        RECT 82.190 66.805 82.580 67.105 ;
        RECT 84.200 66.355 84.370 73.120 ;
        RECT 84.545 71.620 84.865 71.880 ;
        RECT 84.620 69.355 84.790 71.620 ;
        RECT 84.510 69.055 84.900 69.355 ;
        RECT 85.040 67.855 85.210 76.120 ;
        RECT 86.355 75.335 86.525 76.575 ;
        RECT 88.900 75.805 89.290 76.105 ;
        RECT 86.280 75.075 86.600 75.335 ;
        RECT 85.385 74.620 85.705 74.880 ;
        RECT 85.460 70.900 85.630 74.620 ;
        RECT 89.950 74.305 90.340 74.605 ;
        RECT 86.245 73.555 86.635 73.855 ;
        RECT 89.470 73.555 89.860 73.855 ;
        RECT 86.355 72.335 86.525 73.555 ;
        RECT 88.900 72.805 89.290 73.105 ;
        RECT 86.280 72.075 86.600 72.335 ;
        RECT 85.395 70.380 85.695 70.900 ;
        RECT 86.355 70.835 86.525 72.075 ;
        RECT 86.280 70.575 86.600 70.835 ;
        RECT 85.385 70.120 85.705 70.380 ;
        RECT 85.460 69.120 85.630 70.120 ;
        RECT 88.900 69.805 89.290 70.105 ;
        RECT 86.280 68.620 86.600 68.880 ;
        RECT 84.930 67.555 85.320 67.855 ;
        RECT 86.355 67.835 86.525 68.620 ;
        RECT 86.280 67.575 86.600 67.835 ;
        RECT 86.310 67.090 86.570 67.410 ;
        RECT 84.090 66.055 84.480 66.355 ;
        RECT 83.240 65.305 83.630 65.605 ;
        RECT 79.570 63.460 79.890 63.720 ;
        RECT 46.020 63.075 46.340 63.335 ;
        RECT 59.440 63.075 59.760 63.335 ;
        RECT 72.860 63.075 73.180 63.335 ;
        RECT 34.455 60.760 35.495 61.710 ;
        RECT 79.645 59.025 79.815 63.460 ;
        RECT 86.355 63.335 86.525 67.090 ;
        RECT 88.900 66.805 89.290 67.105 ;
        RECT 88.085 65.620 88.405 65.880 ;
        RECT 88.160 63.720 88.330 65.620 ;
        RECT 89.580 64.490 89.750 73.555 ;
        RECT 90.910 73.380 91.080 77.620 ;
        RECT 93.065 76.835 93.235 78.055 ;
        RECT 97.545 77.620 97.865 77.880 ;
        RECT 96.660 77.305 97.050 77.605 ;
        RECT 92.990 76.575 93.310 76.835 ;
        RECT 91.675 76.120 91.995 76.380 ;
        RECT 90.835 73.120 91.155 73.380 ;
        RECT 89.950 71.305 90.340 71.605 ;
        RECT 89.950 68.305 90.340 68.605 ;
        RECT 90.910 66.355 91.080 73.120 ;
        RECT 91.255 71.620 91.575 71.880 ;
        RECT 91.330 69.355 91.500 71.620 ;
        RECT 91.220 69.055 91.610 69.355 ;
        RECT 91.750 67.855 91.920 76.120 ;
        RECT 93.065 75.335 93.235 76.575 ;
        RECT 95.610 75.805 96.000 76.105 ;
        RECT 92.990 75.290 93.310 75.335 ;
        RECT 92.645 75.120 93.310 75.290 ;
        RECT 92.095 74.620 92.415 74.880 ;
        RECT 92.170 70.380 92.340 74.620 ;
        RECT 92.095 70.120 92.415 70.380 ;
        RECT 92.170 68.240 92.340 70.120 ;
        RECT 92.100 67.980 92.420 68.240 ;
        RECT 91.640 67.555 92.030 67.855 ;
        RECT 92.170 67.620 92.340 67.980 ;
        RECT 90.800 66.055 91.190 66.355 ;
        RECT 89.950 65.305 90.340 65.605 ;
        RECT 92.645 64.875 92.815 75.120 ;
        RECT 92.990 75.075 93.310 75.120 ;
        RECT 96.660 74.305 97.050 74.605 ;
        RECT 92.955 73.555 93.345 73.855 ;
        RECT 96.180 73.555 96.570 73.855 ;
        RECT 93.065 72.335 93.235 73.555 ;
        RECT 95.610 72.805 96.000 73.105 ;
        RECT 92.990 72.075 93.310 72.335 ;
        RECT 93.065 70.835 93.235 72.075 ;
        RECT 92.990 70.575 93.310 70.835 ;
        RECT 94.760 70.555 95.150 70.855 ;
        RECT 94.870 69.335 95.040 70.555 ;
        RECT 95.610 69.805 96.000 70.105 ;
        RECT 94.795 69.075 95.115 69.335 ;
        RECT 92.990 68.620 93.310 68.880 ;
        RECT 93.065 67.835 93.235 68.620 ;
        RECT 92.990 67.575 93.310 67.835 ;
        RECT 93.020 67.090 93.280 67.410 ;
        RECT 92.570 64.615 92.890 64.875 ;
        RECT 89.505 64.230 89.825 64.490 ;
        RECT 88.085 63.460 88.405 63.720 ;
        RECT 86.280 63.075 86.600 63.335 ;
        RECT 86.355 59.435 86.525 63.075 ;
        RECT 93.065 59.845 93.235 67.090 ;
        RECT 95.610 66.805 96.000 67.105 ;
        RECT 96.290 63.720 96.460 73.555 ;
        RECT 97.620 73.380 97.790 77.620 ;
        RECT 99.775 76.835 99.945 78.055 ;
        RECT 99.700 76.575 100.020 76.835 ;
        RECT 98.385 76.120 98.705 76.380 ;
        RECT 97.545 73.120 97.865 73.380 ;
        RECT 96.660 71.305 97.050 71.605 ;
        RECT 96.660 68.305 97.050 68.605 ;
        RECT 97.620 66.355 97.790 73.120 ;
        RECT 97.965 71.620 98.285 71.880 ;
        RECT 98.040 69.355 98.210 71.620 ;
        RECT 97.930 69.055 98.320 69.355 ;
        RECT 98.460 67.855 98.630 76.120 ;
        RECT 99.775 75.335 99.945 76.575 ;
        RECT 102.320 75.805 102.710 76.105 ;
        RECT 105.360 76.095 105.660 84.395 ;
        RECT 107.680 83.195 107.980 89.440 ;
        RECT 106.860 82.895 107.980 83.195 ;
        RECT 106.860 77.595 107.160 82.895 ;
        RECT 106.825 77.315 107.195 77.595 ;
        RECT 105.325 75.815 105.695 76.095 ;
        RECT 99.700 75.290 100.020 75.335 ;
        RECT 99.355 75.120 100.020 75.290 ;
        RECT 98.805 74.620 99.125 74.880 ;
        RECT 98.880 70.900 99.050 74.620 ;
        RECT 98.815 70.380 99.115 70.900 ;
        RECT 98.805 70.120 99.125 70.380 ;
        RECT 98.880 69.120 99.050 70.120 ;
        RECT 98.350 67.555 98.740 67.855 ;
        RECT 97.510 66.055 97.900 66.355 ;
        RECT 96.660 65.305 97.050 65.605 ;
        RECT 99.355 64.105 99.525 75.120 ;
        RECT 99.700 75.075 100.020 75.120 ;
        RECT 99.665 73.555 100.055 73.855 ;
        RECT 99.775 72.335 99.945 73.555 ;
        RECT 102.320 72.805 102.710 73.105 ;
        RECT 105.360 73.095 105.660 75.815 ;
        RECT 106.860 74.595 107.160 77.315 ;
        RECT 106.825 74.315 107.195 74.595 ;
        RECT 105.325 72.815 105.695 73.095 ;
        RECT 99.700 72.075 100.020 72.335 ;
        RECT 99.775 70.835 99.945 72.075 ;
        RECT 99.700 70.575 100.020 70.835 ;
        RECT 102.320 69.805 102.710 70.105 ;
        RECT 105.360 70.095 105.660 72.815 ;
        RECT 106.860 71.595 107.160 74.315 ;
        RECT 106.825 71.315 107.195 71.595 ;
        RECT 105.325 69.815 105.695 70.095 ;
        RECT 99.700 68.620 100.020 68.880 ;
        RECT 99.775 67.835 99.945 68.620 ;
        RECT 99.700 67.575 100.020 67.835 ;
        RECT 99.730 67.090 99.990 67.410 ;
        RECT 99.280 63.845 99.600 64.105 ;
        RECT 96.215 63.460 96.535 63.720 ;
        RECT 99.775 60.255 99.945 67.090 ;
        RECT 102.320 66.805 102.710 67.105 ;
        RECT 105.360 67.095 105.660 69.815 ;
        RECT 106.860 68.595 107.160 71.315 ;
        RECT 106.825 68.315 107.195 68.595 ;
        RECT 105.325 66.815 105.695 67.095 ;
        RECT 101.505 65.595 101.825 65.880 ;
        RECT 101.480 65.315 101.850 65.595 ;
        RECT 101.505 65.305 101.825 65.315 ;
        RECT 101.580 65.000 101.750 65.305 ;
        RECT 105.360 61.710 105.660 66.815 ;
        RECT 106.860 65.595 107.160 68.315 ;
        RECT 106.825 65.315 107.195 65.595 ;
        RECT 106.860 63.710 107.160 65.315 ;
        RECT 106.495 62.760 107.535 63.710 ;
        RECT 104.985 60.760 106.025 61.710 ;
        RECT 110.965 60.255 111.245 60.355 ;
        RECT 99.775 60.085 111.245 60.255 ;
        RECT 110.965 59.985 111.245 60.085 ;
        RECT 110.335 59.845 110.615 59.945 ;
        RECT 93.065 59.675 110.615 59.845 ;
        RECT 110.335 59.575 110.615 59.675 ;
        RECT 112.225 59.435 112.505 59.535 ;
        RECT 86.355 59.265 112.505 59.435 ;
        RECT 112.225 59.165 112.505 59.265 ;
        RECT 111.595 59.025 111.875 59.125 ;
        RECT 79.645 58.855 111.875 59.025 ;
        RECT 111.595 58.755 111.875 58.855 ;
      LAYER met3 ;
        RECT 14.990 224.750 15.370 225.070 ;
        RECT 17.750 224.750 18.130 225.070 ;
        RECT 20.510 224.750 20.890 225.070 ;
        RECT 23.270 224.750 23.650 225.070 ;
        RECT 26.030 224.750 26.410 225.070 ;
        RECT 28.790 224.750 29.170 225.070 ;
        RECT 31.550 224.750 31.930 225.070 ;
        RECT 34.310 224.750 34.690 225.070 ;
        RECT 37.070 224.750 37.450 225.070 ;
        RECT 39.830 224.750 40.210 225.070 ;
        RECT 42.590 224.750 42.970 225.070 ;
        RECT 45.350 224.750 45.730 225.070 ;
        RECT 48.110 224.750 48.490 225.070 ;
        RECT 50.870 224.750 51.250 225.070 ;
        RECT 53.630 224.750 54.010 225.070 ;
        RECT 56.390 224.750 56.770 225.070 ;
        RECT 59.150 224.750 59.530 225.070 ;
        RECT 61.910 224.750 62.290 225.070 ;
        RECT 64.670 224.750 65.050 225.070 ;
        RECT 67.430 224.750 67.810 225.070 ;
        RECT 70.190 224.750 70.570 225.070 ;
        RECT 72.950 224.750 73.330 225.070 ;
        RECT 75.710 224.750 76.090 225.070 ;
        RECT 78.470 224.750 78.850 225.070 ;
        RECT 103.310 224.750 103.690 225.070 ;
        RECT 106.070 224.750 106.450 225.070 ;
        RECT 108.830 224.750 109.210 225.070 ;
        RECT 111.590 224.750 111.970 225.070 ;
        RECT 114.350 224.750 114.730 225.070 ;
        RECT 117.110 224.750 117.490 225.070 ;
        RECT 119.870 224.760 120.250 225.080 ;
        RECT 15.030 208.880 15.330 224.750 ;
        RECT 17.790 209.880 18.090 224.750 ;
        RECT 20.550 210.880 20.850 224.750 ;
        RECT 23.310 211.880 23.610 224.750 ;
        RECT 26.070 211.880 26.370 224.750 ;
        RECT 23.310 211.580 24.445 211.880 ;
        RECT 20.550 210.580 22.945 210.880 ;
        RECT 17.790 209.580 21.445 209.880 ;
        RECT 15.030 208.580 19.945 208.880 ;
        RECT 19.645 203.185 19.945 208.580 ;
        RECT 21.145 203.185 21.445 209.580 ;
        RECT 22.645 203.185 22.945 210.580 ;
        RECT 24.145 203.185 24.445 211.580 ;
        RECT 25.645 211.580 26.370 211.880 ;
        RECT 25.645 203.185 25.945 211.580 ;
        RECT 28.830 210.880 29.130 224.750 ;
        RECT 27.145 210.580 29.130 210.880 ;
        RECT 27.145 203.185 27.445 210.580 ;
        RECT 31.590 209.880 31.890 224.750 ;
        RECT 28.645 209.580 31.890 209.880 ;
        RECT 28.645 203.185 28.945 209.580 ;
        RECT 34.350 208.880 34.650 224.750 ;
        RECT 30.145 208.580 34.650 208.880 ;
        RECT 37.110 208.880 37.410 224.750 ;
        RECT 39.870 209.880 40.170 224.750 ;
        RECT 42.630 210.880 42.930 224.750 ;
        RECT 45.390 211.880 45.690 224.750 ;
        RECT 48.150 211.880 48.450 224.750 ;
        RECT 45.390 211.580 46.525 211.880 ;
        RECT 42.630 210.580 45.025 210.880 ;
        RECT 39.870 209.580 43.525 209.880 ;
        RECT 37.110 208.580 42.025 208.880 ;
        RECT 30.145 203.185 30.445 208.580 ;
        RECT 41.725 203.185 42.025 208.580 ;
        RECT 43.225 203.185 43.525 209.580 ;
        RECT 44.725 203.185 45.025 210.580 ;
        RECT 46.225 203.185 46.525 211.580 ;
        RECT 47.725 211.580 48.450 211.880 ;
        RECT 47.725 203.185 48.025 211.580 ;
        RECT 50.910 210.880 51.210 224.750 ;
        RECT 49.225 210.580 51.210 210.880 ;
        RECT 49.225 203.185 49.525 210.580 ;
        RECT 53.670 209.880 53.970 224.750 ;
        RECT 50.725 209.580 53.970 209.880 ;
        RECT 50.725 203.185 51.025 209.580 ;
        RECT 56.430 208.880 56.730 224.750 ;
        RECT 52.225 208.580 56.730 208.880 ;
        RECT 59.190 208.880 59.490 224.750 ;
        RECT 61.950 209.880 62.250 224.750 ;
        RECT 64.710 210.880 65.010 224.750 ;
        RECT 67.470 211.880 67.770 224.750 ;
        RECT 70.230 211.880 70.530 224.750 ;
        RECT 67.470 211.580 68.605 211.880 ;
        RECT 64.710 210.580 67.105 210.880 ;
        RECT 61.950 209.580 65.605 209.880 ;
        RECT 59.190 208.580 64.105 208.880 ;
        RECT 52.225 203.185 52.525 208.580 ;
        RECT 63.805 203.185 64.105 208.580 ;
        RECT 65.305 203.185 65.605 209.580 ;
        RECT 66.805 203.185 67.105 210.580 ;
        RECT 68.305 203.185 68.605 211.580 ;
        RECT 69.805 211.580 70.530 211.880 ;
        RECT 69.805 203.185 70.105 211.580 ;
        RECT 72.990 210.880 73.290 224.750 ;
        RECT 71.305 210.580 73.290 210.880 ;
        RECT 71.305 203.185 71.605 210.580 ;
        RECT 75.750 209.880 76.050 224.750 ;
        RECT 72.805 209.580 76.050 209.880 ;
        RECT 72.805 203.185 73.105 209.580 ;
        RECT 78.510 208.880 78.810 224.750 ;
        RECT 74.305 208.580 78.810 208.880 ;
        RECT 103.350 208.875 103.650 224.750 ;
        RECT 106.110 209.875 106.410 224.750 ;
        RECT 108.870 210.875 109.170 224.750 ;
        RECT 111.630 211.860 111.930 224.750 ;
        RECT 114.390 211.875 114.690 224.750 ;
        RECT 111.630 211.560 112.525 211.860 ;
        RECT 108.870 210.575 111.025 210.875 ;
        RECT 106.110 209.575 109.525 209.875 ;
        RECT 74.305 203.185 74.605 208.580 ;
        RECT 103.350 208.575 108.025 208.875 ;
        RECT 107.725 207.125 108.025 208.575 ;
        RECT 109.225 207.125 109.525 209.575 ;
        RECT 110.725 207.125 111.025 210.575 ;
        RECT 112.225 207.125 112.525 211.560 ;
        RECT 113.725 211.575 114.690 211.875 ;
        RECT 113.725 207.125 114.025 211.575 ;
        RECT 117.150 210.875 117.450 224.750 ;
        RECT 115.225 210.575 117.450 210.875 ;
        RECT 115.225 207.125 115.525 210.575 ;
        RECT 119.910 209.875 120.210 224.760 ;
        RECT 122.630 224.750 123.010 225.070 ;
        RECT 116.725 209.575 120.210 209.875 ;
        RECT 116.725 207.125 117.025 209.575 ;
        RECT 122.670 208.875 122.970 224.750 ;
        RECT 118.225 208.575 122.970 208.875 ;
        RECT 118.225 207.125 118.525 208.575 ;
        RECT 107.710 206.795 108.040 207.125 ;
        RECT 109.210 206.795 109.540 207.125 ;
        RECT 110.710 206.795 111.040 207.125 ;
        RECT 112.210 206.795 112.540 207.125 ;
        RECT 113.710 206.795 114.040 207.125 ;
        RECT 115.210 206.795 115.540 207.125 ;
        RECT 116.710 206.795 117.040 207.125 ;
        RECT 118.210 206.795 118.540 207.125 ;
        RECT 98.500 204.420 99.500 204.450 ;
        RECT 106.395 204.420 107.395 204.445 ;
        RECT 118.920 204.420 119.920 204.445 ;
        RECT 98.500 203.420 120.695 204.420 ;
        RECT 98.500 203.400 99.500 203.420 ;
        RECT 106.395 203.395 107.395 203.420 ;
        RECT 118.920 203.395 119.920 203.420 ;
        RECT 19.630 202.855 19.960 203.185 ;
        RECT 21.130 202.855 21.460 203.185 ;
        RECT 22.630 202.855 22.960 203.185 ;
        RECT 24.130 202.855 24.460 203.185 ;
        RECT 25.630 202.855 25.960 203.185 ;
        RECT 27.130 202.855 27.460 203.185 ;
        RECT 28.630 202.855 28.960 203.185 ;
        RECT 30.130 202.855 30.460 203.185 ;
        RECT 41.710 202.855 42.040 203.185 ;
        RECT 43.210 202.855 43.540 203.185 ;
        RECT 44.710 202.855 45.040 203.185 ;
        RECT 46.210 202.855 46.540 203.185 ;
        RECT 47.710 202.855 48.040 203.185 ;
        RECT 49.210 202.855 49.540 203.185 ;
        RECT 50.710 202.855 51.040 203.185 ;
        RECT 52.210 202.855 52.540 203.185 ;
        RECT 63.790 202.855 64.120 203.185 ;
        RECT 65.290 202.855 65.620 203.185 ;
        RECT 66.790 202.855 67.120 203.185 ;
        RECT 68.290 202.855 68.620 203.185 ;
        RECT 69.790 202.855 70.120 203.185 ;
        RECT 71.290 202.855 71.620 203.185 ;
        RECT 72.790 202.855 73.120 203.185 ;
        RECT 74.290 202.855 74.620 203.185 ;
        RECT 101.500 202.420 102.500 202.450 ;
        RECT 105.145 202.420 106.145 202.445 ;
        RECT 120.170 202.420 121.170 202.445 ;
        RECT 101.500 201.420 121.170 202.420 ;
        RECT 101.500 201.400 102.500 201.420 ;
        RECT 105.145 201.395 106.145 201.420 ;
        RECT 120.170 201.395 121.170 201.420 ;
        RECT 32.500 200.420 33.500 200.450 ;
        RECT 65.500 200.420 66.500 200.450 ;
        RECT 104.500 200.420 105.500 200.450 ;
        RECT 106.395 200.420 107.395 200.445 ;
        RECT 18.600 199.420 75.240 200.420 ;
        RECT 104.500 199.420 120.695 200.420 ;
        RECT 32.500 199.400 33.500 199.420 ;
        RECT 65.500 199.400 66.500 199.420 ;
        RECT 104.500 199.400 105.500 199.420 ;
        RECT 106.395 199.395 107.395 199.420 ;
        RECT 35.500 198.420 36.500 198.450 ;
        RECT 68.500 198.420 69.500 198.450 ;
        RECT 17.350 197.420 76.490 198.420 ;
        RECT 35.500 197.400 36.500 197.420 ;
        RECT 68.500 197.400 69.500 197.420 ;
        RECT 104.500 192.420 105.500 192.450 ;
        RECT 118.920 192.420 119.920 192.445 ;
        RECT 104.500 191.420 120.695 192.420 ;
        RECT 104.500 191.400 105.500 191.420 ;
        RECT 118.920 191.395 119.920 191.420 ;
        RECT 108.165 189.015 108.495 189.345 ;
        RECT 109.665 189.015 109.995 189.345 ;
        RECT 111.165 189.015 111.495 189.345 ;
        RECT 112.665 189.015 112.995 189.345 ;
        RECT 114.165 189.015 114.495 189.345 ;
        RECT 115.665 189.015 115.995 189.345 ;
        RECT 117.165 189.015 117.495 189.345 ;
        RECT 118.665 189.015 118.995 189.345 ;
        RECT 108.180 185.000 108.480 189.015 ;
        RECT 109.680 186.000 109.980 189.015 ;
        RECT 111.180 187.000 111.480 189.015 ;
        RECT 112.680 187.000 112.980 189.015 ;
        RECT 111.180 186.700 111.885 187.000 ;
        RECT 109.680 185.700 111.255 186.000 ;
        RECT 108.180 184.700 110.625 185.000 ;
        RECT 38.500 160.645 39.500 160.675 ;
        RECT 71.500 160.645 72.500 160.675 ;
        RECT 104.500 160.645 105.500 160.675 ;
        RECT 30.325 159.645 108.305 160.645 ;
        RECT 38.500 159.625 39.500 159.645 ;
        RECT 71.500 159.625 72.500 159.645 ;
        RECT 104.500 159.625 105.500 159.645 ;
        RECT 35.500 158.645 36.500 158.675 ;
        RECT 68.500 158.645 69.500 158.675 ;
        RECT 101.500 158.645 102.500 158.675 ;
        RECT 30.325 157.645 108.305 158.645 ;
        RECT 35.500 157.625 36.500 157.645 ;
        RECT 68.500 157.625 69.500 157.645 ;
        RECT 101.500 157.625 102.500 157.645 ;
        RECT 32.500 156.645 33.500 156.675 ;
        RECT 65.500 156.645 66.500 156.675 ;
        RECT 98.500 156.645 99.500 156.675 ;
        RECT 30.325 155.645 108.305 156.645 ;
        RECT 32.500 155.625 33.500 155.645 ;
        RECT 65.500 155.625 66.500 155.645 ;
        RECT 98.500 155.625 99.500 155.645 ;
        RECT 33.130 154.020 33.460 154.035 ;
        RECT 36.975 154.020 37.305 154.035 ;
        RECT 41.775 154.020 42.125 154.045 ;
        RECT 48.485 154.020 48.835 154.045 ;
        RECT 55.195 154.020 55.545 154.045 ;
        RECT 61.905 154.020 62.255 154.045 ;
        RECT 68.615 154.020 68.965 154.045 ;
        RECT 75.325 154.020 75.675 154.045 ;
        RECT 82.035 154.020 82.385 154.045 ;
        RECT 88.745 154.020 89.095 154.045 ;
        RECT 95.455 154.020 95.805 154.045 ;
        RECT 102.165 154.020 102.515 154.045 ;
        RECT 105.170 154.020 105.500 154.035 ;
        RECT 33.130 153.720 105.500 154.020 ;
        RECT 33.130 153.705 33.460 153.720 ;
        RECT 36.975 153.705 37.305 153.720 ;
        RECT 41.775 153.695 42.125 153.720 ;
        RECT 48.485 153.695 48.835 153.720 ;
        RECT 55.195 153.695 55.545 153.720 ;
        RECT 61.905 153.695 62.255 153.720 ;
        RECT 68.615 153.695 68.965 153.720 ;
        RECT 75.325 153.695 75.675 153.720 ;
        RECT 82.035 153.695 82.385 153.720 ;
        RECT 88.745 153.695 89.095 153.720 ;
        RECT 95.455 153.695 95.805 153.720 ;
        RECT 102.165 153.695 102.515 153.720 ;
        RECT 105.170 153.705 105.500 153.720 ;
        RECT 40.925 153.270 41.275 153.295 ;
        RECT 47.635 153.270 47.985 153.295 ;
        RECT 40.925 152.970 47.985 153.270 ;
        RECT 40.925 152.945 41.275 152.970 ;
        RECT 47.635 152.945 47.985 152.970 ;
        RECT 54.345 153.270 54.695 153.295 ;
        RECT 61.055 153.270 61.405 153.295 ;
        RECT 54.345 152.970 61.405 153.270 ;
        RECT 54.345 152.945 54.695 152.970 ;
        RECT 61.055 152.945 61.405 152.970 ;
        RECT 67.765 153.270 68.115 153.295 ;
        RECT 74.475 153.270 74.825 153.295 ;
        RECT 67.765 152.970 74.825 153.270 ;
        RECT 67.765 152.945 68.115 152.970 ;
        RECT 74.475 152.945 74.825 152.970 ;
        RECT 81.185 153.270 81.535 153.295 ;
        RECT 87.895 153.270 88.245 153.295 ;
        RECT 81.185 152.970 88.245 153.270 ;
        RECT 81.185 152.945 81.535 152.970 ;
        RECT 87.895 152.945 88.245 152.970 ;
        RECT 94.605 153.270 94.955 153.295 ;
        RECT 101.315 153.270 101.665 153.295 ;
        RECT 94.605 152.970 101.665 153.270 ;
        RECT 94.605 152.945 94.955 152.970 ;
        RECT 101.315 152.945 101.665 152.970 ;
        RECT 34.630 152.520 34.960 152.535 ;
        RECT 36.115 152.520 36.465 152.545 ;
        RECT 42.825 152.520 43.175 152.545 ;
        RECT 49.535 152.520 49.885 152.545 ;
        RECT 56.245 152.520 56.595 152.545 ;
        RECT 62.955 152.520 63.305 152.545 ;
        RECT 69.665 152.520 70.015 152.545 ;
        RECT 76.375 152.520 76.725 152.545 ;
        RECT 83.085 152.520 83.435 152.545 ;
        RECT 89.795 152.520 90.145 152.545 ;
        RECT 96.505 152.520 96.855 152.545 ;
        RECT 103.670 152.520 104.000 152.535 ;
        RECT 34.630 152.220 104.000 152.520 ;
        RECT 34.630 152.205 34.960 152.220 ;
        RECT 36.115 152.195 36.465 152.220 ;
        RECT 42.825 152.195 43.175 152.220 ;
        RECT 49.535 152.195 49.885 152.220 ;
        RECT 56.245 152.195 56.595 152.220 ;
        RECT 62.955 152.195 63.305 152.220 ;
        RECT 69.665 152.195 70.015 152.220 ;
        RECT 76.375 152.195 76.725 152.220 ;
        RECT 83.085 152.195 83.435 152.220 ;
        RECT 89.795 152.195 90.145 152.220 ;
        RECT 96.505 152.195 96.855 152.220 ;
        RECT 103.670 152.205 104.000 152.220 ;
        RECT 40.085 151.770 40.435 151.795 ;
        RECT 46.795 151.770 47.145 151.795 ;
        RECT 40.085 151.470 47.145 151.770 ;
        RECT 40.085 151.445 40.435 151.470 ;
        RECT 46.795 151.445 47.145 151.470 ;
        RECT 53.505 151.770 53.855 151.795 ;
        RECT 60.215 151.770 60.565 151.795 ;
        RECT 53.505 151.470 60.565 151.770 ;
        RECT 53.505 151.445 53.855 151.470 ;
        RECT 60.215 151.445 60.565 151.470 ;
        RECT 66.925 151.770 67.275 151.795 ;
        RECT 73.635 151.770 73.985 151.795 ;
        RECT 66.925 151.470 73.985 151.770 ;
        RECT 66.925 151.445 67.275 151.470 ;
        RECT 73.635 151.445 73.985 151.470 ;
        RECT 80.345 151.770 80.695 151.795 ;
        RECT 87.055 151.770 87.405 151.795 ;
        RECT 80.345 151.470 87.405 151.770 ;
        RECT 80.345 151.445 80.695 151.470 ;
        RECT 87.055 151.445 87.405 151.470 ;
        RECT 93.765 151.770 94.115 151.795 ;
        RECT 100.475 151.770 100.825 151.795 ;
        RECT 93.765 151.470 100.825 151.770 ;
        RECT 93.765 151.445 94.115 151.470 ;
        RECT 100.475 151.445 100.825 151.470 ;
        RECT 33.130 151.020 33.460 151.035 ;
        RECT 41.775 151.020 42.125 151.045 ;
        RECT 48.485 151.020 48.835 151.045 ;
        RECT 55.195 151.020 55.545 151.045 ;
        RECT 61.905 151.020 62.255 151.045 ;
        RECT 68.615 151.020 68.965 151.045 ;
        RECT 75.325 151.020 75.675 151.045 ;
        RECT 82.035 151.020 82.385 151.045 ;
        RECT 88.745 151.020 89.095 151.045 ;
        RECT 95.455 151.020 95.805 151.045 ;
        RECT 102.165 151.020 102.515 151.045 ;
        RECT 105.170 151.020 105.500 151.035 ;
        RECT 33.130 150.720 105.500 151.020 ;
        RECT 33.130 150.705 33.460 150.720 ;
        RECT 41.775 150.695 42.125 150.720 ;
        RECT 48.485 150.695 48.835 150.720 ;
        RECT 55.195 150.695 55.545 150.720 ;
        RECT 61.905 150.695 62.255 150.720 ;
        RECT 68.615 150.695 68.965 150.720 ;
        RECT 75.325 150.695 75.675 150.720 ;
        RECT 82.035 150.695 82.385 150.720 ;
        RECT 88.745 150.695 89.095 150.720 ;
        RECT 95.455 150.695 95.805 150.720 ;
        RECT 102.165 150.695 102.515 150.720 ;
        RECT 105.170 150.705 105.500 150.720 ;
        RECT 40.505 150.270 40.855 150.295 ;
        RECT 47.215 150.270 47.565 150.295 ;
        RECT 40.505 149.970 47.565 150.270 ;
        RECT 40.505 149.945 40.855 149.970 ;
        RECT 47.215 149.945 47.565 149.970 ;
        RECT 53.925 150.270 54.275 150.295 ;
        RECT 60.635 150.270 60.985 150.295 ;
        RECT 53.925 149.970 60.985 150.270 ;
        RECT 53.925 149.945 54.275 149.970 ;
        RECT 60.635 149.945 60.985 149.970 ;
        RECT 67.345 150.270 67.695 150.295 ;
        RECT 74.055 150.270 74.405 150.295 ;
        RECT 67.345 149.970 74.405 150.270 ;
        RECT 67.345 149.945 67.695 149.970 ;
        RECT 74.055 149.945 74.405 149.970 ;
        RECT 80.765 150.270 81.115 150.295 ;
        RECT 87.475 150.270 87.825 150.295 ;
        RECT 80.765 149.970 87.825 150.270 ;
        RECT 80.765 149.945 81.115 149.970 ;
        RECT 87.475 149.945 87.825 149.970 ;
        RECT 94.185 150.270 94.535 150.295 ;
        RECT 100.895 150.270 101.245 150.295 ;
        RECT 94.185 149.970 101.245 150.270 ;
        RECT 94.185 149.945 94.535 149.970 ;
        RECT 100.895 149.945 101.245 149.970 ;
        RECT 34.630 149.520 34.960 149.535 ;
        RECT 36.115 149.520 36.465 149.545 ;
        RECT 42.825 149.520 43.175 149.545 ;
        RECT 49.535 149.520 49.885 149.545 ;
        RECT 56.245 149.520 56.595 149.545 ;
        RECT 62.955 149.520 63.305 149.545 ;
        RECT 69.665 149.520 70.015 149.545 ;
        RECT 76.375 149.520 76.725 149.545 ;
        RECT 83.085 149.520 83.435 149.545 ;
        RECT 89.795 149.520 90.145 149.545 ;
        RECT 96.505 149.520 96.855 149.545 ;
        RECT 103.670 149.520 104.000 149.535 ;
        RECT 34.630 149.220 104.000 149.520 ;
        RECT 34.630 149.205 34.960 149.220 ;
        RECT 36.115 149.195 36.465 149.220 ;
        RECT 42.825 149.195 43.175 149.220 ;
        RECT 49.535 149.195 49.885 149.220 ;
        RECT 56.245 149.195 56.595 149.220 ;
        RECT 62.955 149.195 63.305 149.220 ;
        RECT 69.665 149.195 70.015 149.220 ;
        RECT 76.375 149.195 76.725 149.220 ;
        RECT 83.085 149.195 83.435 149.220 ;
        RECT 89.795 149.195 90.145 149.220 ;
        RECT 96.505 149.195 96.855 149.220 ;
        RECT 103.670 149.205 104.000 149.220 ;
        RECT 39.665 148.770 40.015 148.795 ;
        RECT 43.675 148.770 44.025 148.795 ;
        RECT 39.665 148.470 44.025 148.770 ;
        RECT 39.665 148.445 40.015 148.470 ;
        RECT 43.675 148.445 44.025 148.470 ;
        RECT 53.085 148.770 53.435 148.795 ;
        RECT 57.095 148.770 57.445 148.795 ;
        RECT 53.085 148.470 57.445 148.770 ;
        RECT 53.085 148.445 53.435 148.470 ;
        RECT 57.095 148.445 57.445 148.470 ;
        RECT 66.505 148.770 66.855 148.795 ;
        RECT 70.515 148.770 70.865 148.795 ;
        RECT 66.505 148.470 70.865 148.770 ;
        RECT 66.505 148.445 66.855 148.470 ;
        RECT 70.515 148.445 70.865 148.470 ;
        RECT 79.925 148.770 80.275 148.795 ;
        RECT 83.935 148.770 84.285 148.795 ;
        RECT 79.925 148.470 84.285 148.770 ;
        RECT 79.925 148.445 80.275 148.470 ;
        RECT 83.935 148.445 84.285 148.470 ;
        RECT 93.345 148.770 93.695 148.795 ;
        RECT 97.355 148.770 97.705 148.795 ;
        RECT 93.345 148.470 97.705 148.770 ;
        RECT 93.345 148.445 93.695 148.470 ;
        RECT 97.355 148.445 97.705 148.470 ;
        RECT 33.130 148.020 33.460 148.035 ;
        RECT 41.775 148.020 42.125 148.045 ;
        RECT 48.485 148.020 48.835 148.045 ;
        RECT 55.195 148.020 55.545 148.045 ;
        RECT 61.905 148.020 62.255 148.045 ;
        RECT 68.615 148.020 68.965 148.045 ;
        RECT 75.325 148.020 75.675 148.045 ;
        RECT 82.035 148.020 82.385 148.045 ;
        RECT 88.745 148.020 89.095 148.045 ;
        RECT 95.455 148.020 95.805 148.045 ;
        RECT 102.165 148.020 102.515 148.045 ;
        RECT 105.170 148.020 105.500 148.035 ;
        RECT 33.130 147.720 105.500 148.020 ;
        RECT 33.130 147.705 33.460 147.720 ;
        RECT 41.775 147.695 42.125 147.720 ;
        RECT 48.485 147.695 48.835 147.720 ;
        RECT 55.195 147.695 55.545 147.720 ;
        RECT 61.905 147.695 62.255 147.720 ;
        RECT 68.615 147.695 68.965 147.720 ;
        RECT 75.325 147.695 75.675 147.720 ;
        RECT 82.035 147.695 82.385 147.720 ;
        RECT 88.745 147.695 89.095 147.720 ;
        RECT 95.455 147.695 95.805 147.720 ;
        RECT 102.165 147.695 102.515 147.720 ;
        RECT 105.170 147.705 105.500 147.720 ;
        RECT 34.630 146.520 34.960 146.535 ;
        RECT 36.115 146.520 36.465 146.545 ;
        RECT 42.825 146.520 43.175 146.545 ;
        RECT 49.535 146.520 49.885 146.545 ;
        RECT 56.245 146.520 56.595 146.545 ;
        RECT 62.955 146.520 63.305 146.545 ;
        RECT 69.665 146.520 70.015 146.545 ;
        RECT 76.375 146.520 76.725 146.545 ;
        RECT 83.085 146.520 83.435 146.545 ;
        RECT 89.795 146.520 90.145 146.545 ;
        RECT 96.505 146.520 96.855 146.545 ;
        RECT 103.670 146.520 104.000 146.535 ;
        RECT 34.630 146.220 104.000 146.520 ;
        RECT 34.630 146.205 34.960 146.220 ;
        RECT 36.115 146.195 36.465 146.220 ;
        RECT 42.825 146.195 43.175 146.220 ;
        RECT 49.535 146.195 49.885 146.220 ;
        RECT 56.245 146.195 56.595 146.220 ;
        RECT 62.955 146.195 63.305 146.220 ;
        RECT 69.665 146.195 70.015 146.220 ;
        RECT 76.375 146.195 76.725 146.220 ;
        RECT 83.085 146.195 83.435 146.220 ;
        RECT 89.795 146.195 90.145 146.220 ;
        RECT 96.505 146.195 96.855 146.220 ;
        RECT 103.670 146.205 104.000 146.220 ;
        RECT 38.770 145.770 39.120 145.795 ;
        RECT 42.255 145.770 42.605 145.795 ;
        RECT 45.480 145.770 45.830 145.795 ;
        RECT 48.965 145.770 49.315 145.795 ;
        RECT 52.190 145.770 52.540 145.795 ;
        RECT 55.675 145.770 56.025 145.795 ;
        RECT 58.900 145.770 59.250 145.795 ;
        RECT 62.385 145.770 62.735 145.795 ;
        RECT 65.610 145.770 65.960 145.795 ;
        RECT 69.095 145.770 69.445 145.795 ;
        RECT 72.320 145.770 72.670 145.795 ;
        RECT 75.805 145.770 76.155 145.795 ;
        RECT 79.030 145.770 79.380 145.795 ;
        RECT 82.515 145.770 82.865 145.795 ;
        RECT 85.740 145.770 86.090 145.795 ;
        RECT 89.225 145.770 89.575 145.795 ;
        RECT 92.450 145.770 92.800 145.795 ;
        RECT 95.935 145.770 96.285 145.795 ;
        RECT 99.160 145.770 99.510 145.795 ;
        RECT 102.645 145.770 102.995 145.795 ;
        RECT 38.275 145.470 42.605 145.770 ;
        RECT 44.985 145.470 49.315 145.770 ;
        RECT 51.695 145.470 56.025 145.770 ;
        RECT 58.405 145.470 62.735 145.770 ;
        RECT 65.115 145.470 69.445 145.770 ;
        RECT 71.825 145.470 76.155 145.770 ;
        RECT 78.535 145.470 82.865 145.770 ;
        RECT 85.245 145.470 89.575 145.770 ;
        RECT 91.955 145.470 96.285 145.770 ;
        RECT 98.665 145.470 102.995 145.770 ;
        RECT 38.770 145.445 39.120 145.470 ;
        RECT 42.255 145.445 42.605 145.470 ;
        RECT 45.480 145.445 45.830 145.470 ;
        RECT 48.965 145.445 49.315 145.470 ;
        RECT 52.190 145.445 52.540 145.470 ;
        RECT 55.675 145.445 56.025 145.470 ;
        RECT 58.900 145.445 59.250 145.470 ;
        RECT 62.385 145.445 62.735 145.470 ;
        RECT 65.610 145.445 65.960 145.470 ;
        RECT 69.095 145.445 69.445 145.470 ;
        RECT 72.320 145.445 72.670 145.470 ;
        RECT 75.805 145.445 76.155 145.470 ;
        RECT 79.030 145.445 79.380 145.470 ;
        RECT 82.515 145.445 82.865 145.470 ;
        RECT 85.740 145.445 86.090 145.470 ;
        RECT 89.225 145.445 89.575 145.470 ;
        RECT 92.450 145.445 92.800 145.470 ;
        RECT 95.935 145.445 96.285 145.470 ;
        RECT 99.160 145.445 99.510 145.470 ;
        RECT 102.645 145.445 102.995 145.470 ;
        RECT 33.130 145.020 33.460 145.035 ;
        RECT 41.775 145.020 42.125 145.045 ;
        RECT 48.485 145.020 48.835 145.045 ;
        RECT 55.195 145.020 55.545 145.045 ;
        RECT 61.905 145.020 62.255 145.045 ;
        RECT 68.615 145.020 68.965 145.045 ;
        RECT 75.325 145.020 75.675 145.045 ;
        RECT 82.035 145.020 82.385 145.045 ;
        RECT 88.745 145.020 89.095 145.045 ;
        RECT 95.455 145.020 95.805 145.045 ;
        RECT 102.165 145.020 102.515 145.045 ;
        RECT 105.170 145.020 105.500 145.035 ;
        RECT 33.130 144.720 105.500 145.020 ;
        RECT 33.130 144.705 33.460 144.720 ;
        RECT 41.775 144.695 42.125 144.720 ;
        RECT 48.485 144.695 48.835 144.720 ;
        RECT 55.195 144.695 55.545 144.720 ;
        RECT 61.905 144.695 62.255 144.720 ;
        RECT 68.615 144.695 68.965 144.720 ;
        RECT 75.325 144.695 75.675 144.720 ;
        RECT 82.035 144.695 82.385 144.720 ;
        RECT 88.745 144.695 89.095 144.720 ;
        RECT 95.455 144.695 95.805 144.720 ;
        RECT 102.165 144.695 102.515 144.720 ;
        RECT 105.170 144.705 105.500 144.720 ;
        RECT 34.630 143.520 34.960 143.535 ;
        RECT 36.115 143.520 36.465 143.545 ;
        RECT 42.825 143.520 43.175 143.545 ;
        RECT 49.535 143.520 49.885 143.545 ;
        RECT 56.245 143.520 56.595 143.545 ;
        RECT 62.955 143.520 63.305 143.545 ;
        RECT 69.665 143.520 70.015 143.545 ;
        RECT 76.375 143.520 76.725 143.545 ;
        RECT 83.085 143.520 83.435 143.545 ;
        RECT 89.795 143.520 90.145 143.545 ;
        RECT 96.505 143.520 96.855 143.545 ;
        RECT 103.670 143.520 104.000 143.535 ;
        RECT 34.630 143.220 104.000 143.520 ;
        RECT 34.630 143.205 34.960 143.220 ;
        RECT 36.115 143.195 36.465 143.220 ;
        RECT 42.825 143.195 43.175 143.220 ;
        RECT 49.535 143.195 49.885 143.220 ;
        RECT 56.245 143.195 56.595 143.220 ;
        RECT 62.955 143.195 63.305 143.220 ;
        RECT 69.665 143.195 70.015 143.220 ;
        RECT 76.375 143.195 76.725 143.220 ;
        RECT 83.085 143.195 83.435 143.220 ;
        RECT 89.795 143.195 90.145 143.220 ;
        RECT 96.505 143.195 96.855 143.220 ;
        RECT 103.670 143.205 104.000 143.220 ;
        RECT 33.130 142.020 33.460 142.035 ;
        RECT 41.775 142.020 42.125 142.045 ;
        RECT 48.485 142.020 48.835 142.045 ;
        RECT 55.195 142.020 55.545 142.045 ;
        RECT 61.905 142.020 62.255 142.045 ;
        RECT 68.615 142.020 68.965 142.045 ;
        RECT 75.325 142.020 75.675 142.045 ;
        RECT 82.035 142.020 82.385 142.045 ;
        RECT 88.745 142.020 89.095 142.045 ;
        RECT 95.455 142.020 95.805 142.045 ;
        RECT 102.165 142.020 102.515 142.045 ;
        RECT 105.170 142.020 105.500 142.035 ;
        RECT 33.130 141.720 105.500 142.020 ;
        RECT 33.130 141.705 33.460 141.720 ;
        RECT 41.775 141.695 42.125 141.720 ;
        RECT 48.485 141.695 48.835 141.720 ;
        RECT 55.195 141.695 55.545 141.720 ;
        RECT 61.905 141.695 62.255 141.720 ;
        RECT 68.615 141.695 68.965 141.720 ;
        RECT 75.325 141.695 75.675 141.720 ;
        RECT 82.035 141.695 82.385 141.720 ;
        RECT 88.745 141.695 89.095 141.720 ;
        RECT 95.455 141.695 95.805 141.720 ;
        RECT 102.165 141.695 102.515 141.720 ;
        RECT 105.170 141.705 105.500 141.720 ;
        RECT 38.770 141.270 39.120 141.295 ;
        RECT 45.480 141.270 45.830 141.295 ;
        RECT 52.190 141.270 52.540 141.295 ;
        RECT 58.900 141.270 59.250 141.295 ;
        RECT 65.610 141.270 65.960 141.295 ;
        RECT 72.320 141.270 72.670 141.295 ;
        RECT 79.030 141.270 79.380 141.295 ;
        RECT 85.740 141.270 86.090 141.295 ;
        RECT 92.450 141.270 92.800 141.295 ;
        RECT 99.160 141.270 99.510 141.295 ;
        RECT 38.275 140.970 39.615 141.270 ;
        RECT 44.985 140.970 46.325 141.270 ;
        RECT 51.695 140.970 53.035 141.270 ;
        RECT 58.405 140.970 59.745 141.270 ;
        RECT 65.115 140.970 66.455 141.270 ;
        RECT 71.825 140.970 73.165 141.270 ;
        RECT 78.535 140.970 79.875 141.270 ;
        RECT 85.245 140.970 86.585 141.270 ;
        RECT 91.955 140.970 93.295 141.270 ;
        RECT 98.665 140.970 100.005 141.270 ;
        RECT 38.770 140.945 39.120 140.970 ;
        RECT 45.480 140.945 45.830 140.970 ;
        RECT 52.190 140.945 52.540 140.970 ;
        RECT 58.900 140.945 59.250 140.970 ;
        RECT 65.610 140.945 65.960 140.970 ;
        RECT 72.320 140.945 72.670 140.970 ;
        RECT 79.030 140.945 79.380 140.970 ;
        RECT 85.740 140.945 86.090 140.970 ;
        RECT 92.450 140.945 92.800 140.970 ;
        RECT 99.160 140.945 99.510 140.970 ;
        RECT 38.500 138.645 39.500 138.675 ;
        RECT 71.500 138.645 72.500 138.675 ;
        RECT 104.500 138.645 105.500 138.675 ;
        RECT 30.325 137.645 108.305 138.645 ;
        RECT 38.500 137.625 39.500 137.645 ;
        RECT 71.500 137.625 72.500 137.645 ;
        RECT 104.500 137.625 105.500 137.645 ;
        RECT 35.500 136.645 36.500 136.675 ;
        RECT 68.500 136.645 69.500 136.675 ;
        RECT 101.500 136.645 102.500 136.675 ;
        RECT 30.325 135.645 108.305 136.645 ;
        RECT 35.500 135.625 36.500 135.645 ;
        RECT 68.500 135.625 69.500 135.645 ;
        RECT 101.500 135.625 102.500 135.645 ;
        RECT 59.785 133.290 60.115 133.620 ;
        RECT 61.165 133.290 61.495 133.620 ;
        RECT 62.545 133.290 62.875 133.620 ;
        RECT 63.925 133.290 64.255 133.620 ;
        RECT 65.305 133.290 65.635 133.620 ;
        RECT 66.685 133.290 67.015 133.620 ;
        RECT 68.065 133.290 68.395 133.620 ;
        RECT 69.445 133.290 69.775 133.620 ;
        RECT 70.825 133.290 71.155 133.620 ;
        RECT 72.205 133.290 72.535 133.620 ;
        RECT 73.585 133.290 73.915 133.620 ;
        RECT 74.965 133.290 75.295 133.620 ;
        RECT 76.345 133.290 76.675 133.620 ;
        RECT 77.725 133.290 78.055 133.620 ;
        RECT 79.105 133.290 79.435 133.620 ;
        RECT 80.485 133.290 80.815 133.620 ;
        RECT 59.800 131.945 60.100 133.290 ;
        RECT 61.180 131.945 61.480 133.290 ;
        RECT 62.560 131.945 62.860 133.290 ;
        RECT 63.940 131.945 64.240 133.290 ;
        RECT 65.320 131.945 65.620 133.290 ;
        RECT 66.700 131.945 67.000 133.290 ;
        RECT 68.080 131.945 68.380 133.290 ;
        RECT 69.460 131.945 69.760 133.290 ;
        RECT 70.840 131.945 71.140 133.290 ;
        RECT 72.220 131.945 72.520 133.290 ;
        RECT 73.600 131.945 73.900 133.290 ;
        RECT 74.980 131.945 75.280 133.290 ;
        RECT 76.360 131.945 76.660 133.290 ;
        RECT 77.740 131.945 78.040 133.290 ;
        RECT 79.120 131.945 79.420 133.290 ;
        RECT 80.500 131.945 80.800 133.290 ;
        RECT 59.775 131.615 60.125 131.945 ;
        RECT 61.155 131.615 61.505 131.945 ;
        RECT 62.535 131.615 62.885 131.945 ;
        RECT 63.915 131.615 64.265 131.945 ;
        RECT 65.295 131.615 65.645 131.945 ;
        RECT 66.675 131.615 67.025 131.945 ;
        RECT 68.055 131.615 68.405 131.945 ;
        RECT 69.435 131.615 69.785 131.945 ;
        RECT 70.815 131.615 71.165 131.945 ;
        RECT 72.195 131.615 72.545 131.945 ;
        RECT 73.575 131.615 73.925 131.945 ;
        RECT 74.955 131.615 75.305 131.945 ;
        RECT 76.335 131.615 76.685 131.945 ;
        RECT 77.715 131.615 78.065 131.945 ;
        RECT 79.095 131.615 79.445 131.945 ;
        RECT 80.475 131.615 80.825 131.945 ;
        RECT 59.495 129.625 108.410 130.525 ;
        RECT 79.990 127.045 80.340 127.075 ;
        RECT 59.240 126.645 59.640 127.045 ;
        RECT 60.620 126.645 61.020 127.045 ;
        RECT 62.000 126.645 62.400 127.045 ;
        RECT 63.380 126.645 63.780 127.045 ;
        RECT 64.760 126.645 65.160 127.045 ;
        RECT 66.140 126.645 66.540 127.045 ;
        RECT 67.520 126.645 67.920 127.045 ;
        RECT 68.900 126.645 69.300 127.045 ;
        RECT 70.280 126.645 70.680 127.045 ;
        RECT 71.660 126.645 72.060 127.045 ;
        RECT 73.040 126.645 73.440 127.045 ;
        RECT 74.420 126.645 74.820 127.045 ;
        RECT 75.800 126.645 76.200 127.045 ;
        RECT 77.180 126.645 77.580 127.045 ;
        RECT 78.560 126.645 78.960 127.045 ;
        RECT 79.940 126.645 80.340 127.045 ;
        RECT 59.265 116.790 59.615 126.645 ;
        RECT 60.645 117.440 60.995 126.645 ;
        RECT 62.025 118.090 62.375 126.645 ;
        RECT 63.405 118.740 63.755 126.645 ;
        RECT 64.785 119.390 65.135 126.645 ;
        RECT 66.165 120.040 66.515 126.645 ;
        RECT 67.545 120.690 67.895 126.645 ;
        RECT 68.925 121.340 69.275 126.645 ;
        RECT 70.305 121.990 70.655 126.645 ;
        RECT 71.685 122.640 72.035 126.645 ;
        RECT 73.065 123.290 73.415 126.645 ;
        RECT 74.445 123.940 74.795 126.645 ;
        RECT 75.825 124.590 76.175 126.645 ;
        RECT 77.205 125.240 77.555 126.645 ;
        RECT 78.585 125.890 78.935 126.645 ;
        RECT 79.965 126.565 80.340 126.645 ;
        RECT 79.965 126.215 82.395 126.565 ;
        RECT 78.585 125.540 81.565 125.890 ;
        RECT 77.205 124.890 80.735 125.240 ;
        RECT 75.825 124.240 79.905 124.590 ;
        RECT 74.445 123.590 79.075 123.940 ;
        RECT 73.065 122.940 78.245 123.290 ;
        RECT 71.685 122.290 77.415 122.640 ;
        RECT 77.065 122.045 77.415 122.290 ;
        RECT 77.895 122.045 78.245 122.940 ;
        RECT 78.725 122.045 79.075 123.590 ;
        RECT 79.555 122.045 79.905 124.240 ;
        RECT 80.385 122.045 80.735 124.890 ;
        RECT 81.215 122.045 81.565 125.540 ;
        RECT 70.305 121.640 76.585 121.990 ;
        RECT 68.925 120.990 75.755 121.340 ;
        RECT 67.545 120.340 74.925 120.690 ;
        RECT 66.165 119.690 74.095 120.040 ;
        RECT 64.785 119.040 73.265 119.390 ;
        RECT 63.405 118.390 72.435 118.740 ;
        RECT 62.025 117.740 71.605 118.090 ;
        RECT 60.645 117.090 70.775 117.440 ;
        RECT 59.265 116.440 69.945 116.790 ;
        RECT 69.570 114.215 69.970 114.240 ;
        RECT 69.570 113.865 81.500 114.215 ;
        RECT 69.570 113.840 69.970 113.865 ;
        RECT 55.550 113.190 80.825 113.540 ;
        RECT 68.765 112.540 79.445 112.890 ;
        RECT 67.935 111.890 78.065 112.240 ;
        RECT 67.105 111.240 76.685 111.590 ;
        RECT 66.275 110.590 75.305 110.940 ;
        RECT 65.445 109.940 73.925 110.290 ;
        RECT 64.615 109.290 72.545 109.640 ;
        RECT 63.785 108.640 71.165 108.990 ;
        RECT 62.955 107.990 69.785 108.340 ;
        RECT 62.125 107.340 68.405 107.690 ;
        RECT 56.315 103.115 56.665 107.285 ;
        RECT 57.145 103.790 57.495 107.285 ;
        RECT 57.975 104.440 58.325 107.285 ;
        RECT 58.805 105.090 59.155 107.285 ;
        RECT 59.635 105.740 59.985 107.285 ;
        RECT 60.465 106.390 60.815 107.285 ;
        RECT 61.295 107.040 61.645 107.285 ;
        RECT 61.295 106.690 67.025 107.040 ;
        RECT 60.465 106.040 65.645 106.390 ;
        RECT 59.635 105.390 64.265 105.740 ;
        RECT 58.805 104.740 62.885 105.090 ;
        RECT 57.975 104.090 61.505 104.440 ;
        RECT 57.145 103.440 60.125 103.790 ;
        RECT 56.315 102.765 58.745 103.115 ;
        RECT 58.370 102.685 58.745 102.765 ;
        RECT 59.775 102.685 60.125 103.440 ;
        RECT 61.155 102.685 61.505 104.090 ;
        RECT 62.535 102.685 62.885 104.740 ;
        RECT 63.915 102.685 64.265 105.390 ;
        RECT 65.295 102.685 65.645 106.040 ;
        RECT 66.675 102.685 67.025 106.690 ;
        RECT 68.055 102.685 68.405 107.340 ;
        RECT 69.435 102.685 69.785 107.990 ;
        RECT 70.815 102.685 71.165 108.640 ;
        RECT 72.195 102.685 72.545 109.290 ;
        RECT 73.575 102.685 73.925 109.940 ;
        RECT 74.955 102.685 75.305 110.590 ;
        RECT 76.335 102.685 76.685 111.240 ;
        RECT 77.715 102.685 78.065 111.890 ;
        RECT 79.095 102.685 79.445 112.540 ;
        RECT 80.475 102.685 80.825 113.190 ;
        RECT 58.370 102.285 58.770 102.685 ;
        RECT 59.750 102.285 60.150 102.685 ;
        RECT 61.130 102.285 61.530 102.685 ;
        RECT 62.510 102.285 62.910 102.685 ;
        RECT 63.890 102.285 64.290 102.685 ;
        RECT 65.270 102.285 65.670 102.685 ;
        RECT 66.650 102.285 67.050 102.685 ;
        RECT 68.030 102.285 68.430 102.685 ;
        RECT 69.410 102.285 69.810 102.685 ;
        RECT 70.790 102.285 71.190 102.685 ;
        RECT 72.170 102.285 72.570 102.685 ;
        RECT 73.550 102.285 73.950 102.685 ;
        RECT 74.930 102.285 75.330 102.685 ;
        RECT 76.310 102.285 76.710 102.685 ;
        RECT 77.690 102.285 78.090 102.685 ;
        RECT 79.070 102.285 79.470 102.685 ;
        RECT 80.450 102.285 80.850 102.685 ;
        RECT 81.150 100.250 81.500 113.865 ;
        RECT 82.045 109.490 82.395 126.215 ;
        RECT 82.020 109.090 82.420 109.490 ;
        RECT 59.265 99.900 81.500 100.250 ;
        RECT 59.265 99.600 59.615 99.900 ;
        RECT 62.025 99.600 62.375 99.900 ;
        RECT 64.785 99.600 65.135 99.900 ;
        RECT 67.545 99.600 67.895 99.900 ;
        RECT 70.305 99.600 70.655 99.900 ;
        RECT 73.065 99.600 73.415 99.900 ;
        RECT 75.825 99.600 76.175 99.900 ;
        RECT 78.585 99.600 78.935 99.900 ;
        RECT 57.715 98.910 58.405 99.600 ;
        RECT 59.095 98.910 59.785 99.600 ;
        RECT 60.475 98.910 61.165 99.600 ;
        RECT 61.855 98.910 62.545 99.600 ;
        RECT 63.235 98.910 63.925 99.600 ;
        RECT 64.615 98.910 65.305 99.600 ;
        RECT 65.995 98.910 66.685 99.600 ;
        RECT 67.375 98.910 68.065 99.600 ;
        RECT 68.755 98.910 69.445 99.600 ;
        RECT 70.135 98.910 70.825 99.600 ;
        RECT 71.515 98.910 72.205 99.600 ;
        RECT 72.895 98.910 73.585 99.600 ;
        RECT 74.275 98.910 74.965 99.600 ;
        RECT 75.655 98.910 76.345 99.600 ;
        RECT 77.035 98.910 77.725 99.600 ;
        RECT 78.415 98.910 79.105 99.600 ;
        RECT 79.795 98.910 80.485 99.600 ;
        RECT 57.885 98.610 58.235 98.910 ;
        RECT 60.645 98.610 60.995 98.910 ;
        RECT 63.405 98.610 63.755 98.910 ;
        RECT 66.165 98.610 66.515 98.910 ;
        RECT 68.925 98.610 69.275 98.910 ;
        RECT 71.685 98.610 72.035 98.910 ;
        RECT 74.445 98.610 74.795 98.910 ;
        RECT 77.205 98.610 77.555 98.910 ;
        RECT 79.965 98.610 80.315 98.910 ;
        RECT 82.045 98.610 82.395 109.090 ;
        RECT 57.885 98.260 82.395 98.610 ;
        RECT 57.885 97.395 58.235 97.725 ;
        RECT 59.265 97.395 59.615 97.725 ;
        RECT 60.645 97.395 60.995 97.725 ;
        RECT 62.025 97.395 62.375 97.725 ;
        RECT 63.405 97.395 63.755 97.725 ;
        RECT 64.785 97.395 65.135 97.725 ;
        RECT 66.165 97.395 66.515 97.725 ;
        RECT 67.545 97.395 67.895 97.725 ;
        RECT 68.925 97.395 69.275 97.725 ;
        RECT 70.305 97.395 70.655 97.725 ;
        RECT 71.685 97.395 72.035 97.725 ;
        RECT 73.065 97.395 73.415 97.725 ;
        RECT 74.445 97.395 74.795 97.725 ;
        RECT 75.825 97.395 76.175 97.725 ;
        RECT 77.205 97.395 77.555 97.725 ;
        RECT 78.585 97.395 78.935 97.725 ;
        RECT 79.965 97.395 80.315 97.725 ;
        RECT 57.910 96.060 58.210 97.395 ;
        RECT 59.290 96.060 59.590 97.395 ;
        RECT 60.670 96.060 60.970 97.395 ;
        RECT 62.050 96.060 62.350 97.395 ;
        RECT 63.430 96.060 63.730 97.395 ;
        RECT 64.810 96.060 65.110 97.395 ;
        RECT 66.190 96.060 66.490 97.395 ;
        RECT 67.570 96.060 67.870 97.395 ;
        RECT 68.950 96.060 69.250 97.395 ;
        RECT 70.330 96.060 70.630 97.395 ;
        RECT 71.710 96.060 72.010 97.395 ;
        RECT 73.090 96.060 73.390 97.395 ;
        RECT 74.470 96.060 74.770 97.395 ;
        RECT 75.850 96.060 76.150 97.395 ;
        RECT 77.230 96.060 77.530 97.395 ;
        RECT 78.610 96.060 78.910 97.395 ;
        RECT 79.990 96.060 80.290 97.395 ;
        RECT 57.895 95.730 58.225 96.060 ;
        RECT 59.275 95.730 59.605 96.060 ;
        RECT 60.655 95.730 60.985 96.060 ;
        RECT 62.035 95.730 62.365 96.060 ;
        RECT 63.415 95.730 63.745 96.060 ;
        RECT 64.795 95.730 65.125 96.060 ;
        RECT 66.175 95.730 66.505 96.060 ;
        RECT 67.555 95.730 67.885 96.060 ;
        RECT 68.935 95.730 69.265 96.060 ;
        RECT 70.315 95.730 70.645 96.060 ;
        RECT 71.695 95.730 72.025 96.060 ;
        RECT 73.075 95.730 73.405 96.060 ;
        RECT 74.455 95.730 74.785 96.060 ;
        RECT 75.835 95.730 76.165 96.060 ;
        RECT 77.215 95.730 77.545 96.060 ;
        RECT 78.595 95.730 78.925 96.060 ;
        RECT 79.975 95.730 80.305 96.060 ;
        RECT 38.500 93.735 39.500 93.765 ;
        RECT 71.500 93.735 72.500 93.765 ;
        RECT 104.500 93.735 105.500 93.765 ;
        RECT 30.325 92.735 108.305 93.735 ;
        RECT 38.500 92.715 39.500 92.735 ;
        RECT 71.500 92.715 72.500 92.735 ;
        RECT 104.500 92.715 105.500 92.735 ;
        RECT 35.500 91.735 36.500 91.765 ;
        RECT 68.500 91.735 69.500 91.765 ;
        RECT 101.500 91.735 102.500 91.765 ;
        RECT 30.325 90.735 108.305 91.735 ;
        RECT 35.500 90.715 36.500 90.735 ;
        RECT 68.500 90.715 69.500 90.735 ;
        RECT 101.500 90.715 102.500 90.735 ;
        RECT 39.295 78.355 39.645 78.380 ;
        RECT 46.005 78.355 46.355 78.380 ;
        RECT 52.715 78.355 53.065 78.380 ;
        RECT 59.425 78.355 59.775 78.380 ;
        RECT 66.135 78.355 66.485 78.380 ;
        RECT 72.845 78.355 73.195 78.380 ;
        RECT 79.555 78.355 79.905 78.380 ;
        RECT 86.265 78.355 86.615 78.380 ;
        RECT 92.975 78.355 93.325 78.380 ;
        RECT 99.685 78.355 100.035 78.380 ;
        RECT 38.800 78.055 40.140 78.355 ;
        RECT 45.510 78.055 46.850 78.355 ;
        RECT 52.220 78.055 53.560 78.355 ;
        RECT 58.930 78.055 60.270 78.355 ;
        RECT 65.640 78.055 66.980 78.355 ;
        RECT 72.350 78.055 73.690 78.355 ;
        RECT 79.060 78.055 80.400 78.355 ;
        RECT 85.770 78.055 87.110 78.355 ;
        RECT 92.480 78.055 93.820 78.355 ;
        RECT 99.190 78.055 100.530 78.355 ;
        RECT 39.295 78.030 39.645 78.055 ;
        RECT 46.005 78.030 46.355 78.055 ;
        RECT 52.715 78.030 53.065 78.055 ;
        RECT 59.425 78.030 59.775 78.055 ;
        RECT 66.135 78.030 66.485 78.055 ;
        RECT 72.845 78.030 73.195 78.055 ;
        RECT 79.555 78.030 79.905 78.055 ;
        RECT 86.265 78.030 86.615 78.055 ;
        RECT 92.975 78.030 93.325 78.055 ;
        RECT 99.685 78.030 100.035 78.055 ;
        RECT 33.305 77.605 33.635 77.620 ;
        RECT 36.290 77.605 36.640 77.630 ;
        RECT 43.000 77.605 43.350 77.630 ;
        RECT 49.710 77.605 50.060 77.630 ;
        RECT 56.420 77.605 56.770 77.630 ;
        RECT 63.130 77.605 63.480 77.630 ;
        RECT 69.840 77.605 70.190 77.630 ;
        RECT 76.550 77.605 76.900 77.630 ;
        RECT 83.260 77.605 83.610 77.630 ;
        RECT 89.970 77.605 90.320 77.630 ;
        RECT 96.680 77.605 97.030 77.630 ;
        RECT 106.845 77.605 107.175 77.620 ;
        RECT 33.305 77.305 107.175 77.605 ;
        RECT 33.305 77.290 33.635 77.305 ;
        RECT 36.290 77.280 36.640 77.305 ;
        RECT 43.000 77.280 43.350 77.305 ;
        RECT 49.710 77.280 50.060 77.305 ;
        RECT 56.420 77.280 56.770 77.305 ;
        RECT 63.130 77.280 63.480 77.305 ;
        RECT 69.840 77.280 70.190 77.305 ;
        RECT 76.550 77.280 76.900 77.305 ;
        RECT 83.260 77.280 83.610 77.305 ;
        RECT 89.970 77.280 90.320 77.305 ;
        RECT 96.680 77.280 97.030 77.305 ;
        RECT 106.845 77.290 107.175 77.305 ;
        RECT 34.805 76.105 35.135 76.120 ;
        RECT 41.950 76.105 42.300 76.130 ;
        RECT 48.660 76.105 49.010 76.130 ;
        RECT 55.370 76.105 55.720 76.130 ;
        RECT 62.080 76.105 62.430 76.130 ;
        RECT 68.790 76.105 69.140 76.130 ;
        RECT 75.500 76.105 75.850 76.130 ;
        RECT 82.210 76.105 82.560 76.130 ;
        RECT 88.920 76.105 89.270 76.130 ;
        RECT 95.630 76.105 95.980 76.130 ;
        RECT 102.340 76.105 102.690 76.130 ;
        RECT 105.345 76.105 105.675 76.120 ;
        RECT 34.805 75.805 105.675 76.105 ;
        RECT 34.805 75.790 35.135 75.805 ;
        RECT 41.950 75.780 42.300 75.805 ;
        RECT 48.660 75.780 49.010 75.805 ;
        RECT 55.370 75.780 55.720 75.805 ;
        RECT 62.080 75.780 62.430 75.805 ;
        RECT 68.790 75.780 69.140 75.805 ;
        RECT 75.500 75.780 75.850 75.805 ;
        RECT 82.210 75.780 82.560 75.805 ;
        RECT 88.920 75.780 89.270 75.805 ;
        RECT 95.630 75.780 95.980 75.805 ;
        RECT 102.340 75.780 102.690 75.805 ;
        RECT 105.345 75.790 105.675 75.805 ;
        RECT 33.305 74.605 33.635 74.620 ;
        RECT 36.290 74.605 36.640 74.630 ;
        RECT 43.000 74.605 43.350 74.630 ;
        RECT 49.710 74.605 50.060 74.630 ;
        RECT 56.420 74.605 56.770 74.630 ;
        RECT 63.130 74.605 63.480 74.630 ;
        RECT 69.840 74.605 70.190 74.630 ;
        RECT 76.550 74.605 76.900 74.630 ;
        RECT 83.260 74.605 83.610 74.630 ;
        RECT 89.970 74.605 90.320 74.630 ;
        RECT 96.680 74.605 97.030 74.630 ;
        RECT 106.845 74.605 107.175 74.620 ;
        RECT 33.305 74.305 107.175 74.605 ;
        RECT 33.305 74.290 33.635 74.305 ;
        RECT 36.290 74.280 36.640 74.305 ;
        RECT 43.000 74.280 43.350 74.305 ;
        RECT 49.710 74.280 50.060 74.305 ;
        RECT 56.420 74.280 56.770 74.305 ;
        RECT 63.130 74.280 63.480 74.305 ;
        RECT 69.840 74.280 70.190 74.305 ;
        RECT 76.550 74.280 76.900 74.305 ;
        RECT 83.260 74.280 83.610 74.305 ;
        RECT 89.970 74.280 90.320 74.305 ;
        RECT 96.680 74.280 97.030 74.305 ;
        RECT 106.845 74.290 107.175 74.305 ;
        RECT 35.810 73.855 36.160 73.880 ;
        RECT 39.295 73.855 39.645 73.880 ;
        RECT 42.520 73.855 42.870 73.880 ;
        RECT 46.005 73.855 46.355 73.880 ;
        RECT 49.230 73.855 49.580 73.880 ;
        RECT 52.715 73.855 53.065 73.880 ;
        RECT 55.940 73.855 56.290 73.880 ;
        RECT 59.425 73.855 59.775 73.880 ;
        RECT 62.650 73.855 63.000 73.880 ;
        RECT 66.135 73.855 66.485 73.880 ;
        RECT 69.360 73.855 69.710 73.880 ;
        RECT 72.845 73.855 73.195 73.880 ;
        RECT 76.070 73.855 76.420 73.880 ;
        RECT 79.555 73.855 79.905 73.880 ;
        RECT 82.780 73.855 83.130 73.880 ;
        RECT 86.265 73.855 86.615 73.880 ;
        RECT 89.490 73.855 89.840 73.880 ;
        RECT 92.975 73.855 93.325 73.880 ;
        RECT 96.200 73.855 96.550 73.880 ;
        RECT 99.685 73.855 100.035 73.880 ;
        RECT 35.810 73.555 40.140 73.855 ;
        RECT 42.520 73.555 46.850 73.855 ;
        RECT 49.230 73.555 53.560 73.855 ;
        RECT 55.940 73.555 60.270 73.855 ;
        RECT 62.650 73.555 66.980 73.855 ;
        RECT 69.360 73.555 73.690 73.855 ;
        RECT 76.070 73.555 80.400 73.855 ;
        RECT 82.780 73.555 87.110 73.855 ;
        RECT 89.490 73.555 93.820 73.855 ;
        RECT 96.200 73.555 100.530 73.855 ;
        RECT 35.810 73.530 36.160 73.555 ;
        RECT 39.295 73.530 39.645 73.555 ;
        RECT 42.520 73.530 42.870 73.555 ;
        RECT 46.005 73.530 46.355 73.555 ;
        RECT 49.230 73.530 49.580 73.555 ;
        RECT 52.715 73.530 53.065 73.555 ;
        RECT 55.940 73.530 56.290 73.555 ;
        RECT 59.425 73.530 59.775 73.555 ;
        RECT 62.650 73.530 63.000 73.555 ;
        RECT 66.135 73.530 66.485 73.555 ;
        RECT 69.360 73.530 69.710 73.555 ;
        RECT 72.845 73.530 73.195 73.555 ;
        RECT 76.070 73.530 76.420 73.555 ;
        RECT 79.555 73.530 79.905 73.555 ;
        RECT 82.780 73.530 83.130 73.555 ;
        RECT 86.265 73.530 86.615 73.555 ;
        RECT 89.490 73.530 89.840 73.555 ;
        RECT 92.975 73.530 93.325 73.555 ;
        RECT 96.200 73.530 96.550 73.555 ;
        RECT 99.685 73.530 100.035 73.555 ;
        RECT 34.805 73.105 35.135 73.120 ;
        RECT 41.950 73.105 42.300 73.130 ;
        RECT 48.660 73.105 49.010 73.130 ;
        RECT 55.370 73.105 55.720 73.130 ;
        RECT 62.080 73.105 62.430 73.130 ;
        RECT 68.790 73.105 69.140 73.130 ;
        RECT 75.500 73.105 75.850 73.130 ;
        RECT 82.210 73.105 82.560 73.130 ;
        RECT 88.920 73.105 89.270 73.130 ;
        RECT 95.630 73.105 95.980 73.130 ;
        RECT 102.340 73.105 102.690 73.130 ;
        RECT 105.345 73.105 105.675 73.120 ;
        RECT 34.805 72.805 105.675 73.105 ;
        RECT 34.805 72.790 35.135 72.805 ;
        RECT 41.950 72.780 42.300 72.805 ;
        RECT 48.660 72.780 49.010 72.805 ;
        RECT 55.370 72.780 55.720 72.805 ;
        RECT 62.080 72.780 62.430 72.805 ;
        RECT 68.790 72.780 69.140 72.805 ;
        RECT 75.500 72.780 75.850 72.805 ;
        RECT 82.210 72.780 82.560 72.805 ;
        RECT 88.920 72.780 89.270 72.805 ;
        RECT 95.630 72.780 95.980 72.805 ;
        RECT 102.340 72.780 102.690 72.805 ;
        RECT 105.345 72.790 105.675 72.805 ;
        RECT 33.305 71.605 33.635 71.620 ;
        RECT 36.290 71.605 36.640 71.630 ;
        RECT 43.000 71.605 43.350 71.630 ;
        RECT 49.710 71.605 50.060 71.630 ;
        RECT 56.420 71.605 56.770 71.630 ;
        RECT 63.130 71.605 63.480 71.630 ;
        RECT 69.840 71.605 70.190 71.630 ;
        RECT 76.550 71.605 76.900 71.630 ;
        RECT 83.260 71.605 83.610 71.630 ;
        RECT 89.970 71.605 90.320 71.630 ;
        RECT 96.680 71.605 97.030 71.630 ;
        RECT 106.845 71.605 107.175 71.620 ;
        RECT 33.305 71.305 107.175 71.605 ;
        RECT 33.305 71.290 33.635 71.305 ;
        RECT 36.290 71.280 36.640 71.305 ;
        RECT 43.000 71.280 43.350 71.305 ;
        RECT 49.710 71.280 50.060 71.305 ;
        RECT 56.420 71.280 56.770 71.305 ;
        RECT 63.130 71.280 63.480 71.305 ;
        RECT 69.840 71.280 70.190 71.305 ;
        RECT 76.550 71.280 76.900 71.305 ;
        RECT 83.260 71.280 83.610 71.305 ;
        RECT 89.970 71.280 90.320 71.305 ;
        RECT 96.680 71.280 97.030 71.305 ;
        RECT 106.845 71.290 107.175 71.305 ;
        RECT 41.100 70.855 41.450 70.880 ;
        RECT 45.110 70.855 45.460 70.880 ;
        RECT 41.100 70.555 45.460 70.855 ;
        RECT 41.100 70.530 41.450 70.555 ;
        RECT 45.110 70.530 45.460 70.555 ;
        RECT 54.520 70.855 54.870 70.880 ;
        RECT 58.530 70.855 58.880 70.880 ;
        RECT 54.520 70.555 58.880 70.855 ;
        RECT 54.520 70.530 54.870 70.555 ;
        RECT 58.530 70.530 58.880 70.555 ;
        RECT 67.940 70.855 68.290 70.880 ;
        RECT 71.950 70.855 72.300 70.880 ;
        RECT 67.940 70.555 72.300 70.855 ;
        RECT 67.940 70.530 68.290 70.555 ;
        RECT 71.950 70.530 72.300 70.555 ;
        RECT 81.360 70.855 81.710 70.880 ;
        RECT 85.370 70.855 85.720 70.880 ;
        RECT 81.360 70.555 85.720 70.855 ;
        RECT 81.360 70.530 81.710 70.555 ;
        RECT 85.370 70.530 85.720 70.555 ;
        RECT 94.780 70.855 95.130 70.880 ;
        RECT 98.790 70.855 99.140 70.880 ;
        RECT 94.780 70.555 99.140 70.855 ;
        RECT 94.780 70.530 95.130 70.555 ;
        RECT 98.790 70.530 99.140 70.555 ;
        RECT 34.805 70.105 35.135 70.120 ;
        RECT 41.950 70.105 42.300 70.130 ;
        RECT 48.660 70.105 49.010 70.130 ;
        RECT 55.370 70.105 55.720 70.130 ;
        RECT 62.080 70.105 62.430 70.130 ;
        RECT 68.790 70.105 69.140 70.130 ;
        RECT 75.500 70.105 75.850 70.130 ;
        RECT 82.210 70.105 82.560 70.130 ;
        RECT 88.920 70.105 89.270 70.130 ;
        RECT 95.630 70.105 95.980 70.130 ;
        RECT 102.340 70.105 102.690 70.130 ;
        RECT 105.345 70.105 105.675 70.120 ;
        RECT 34.805 69.805 105.675 70.105 ;
        RECT 34.805 69.790 35.135 69.805 ;
        RECT 41.950 69.780 42.300 69.805 ;
        RECT 48.660 69.780 49.010 69.805 ;
        RECT 55.370 69.780 55.720 69.805 ;
        RECT 62.080 69.780 62.430 69.805 ;
        RECT 68.790 69.780 69.140 69.805 ;
        RECT 75.500 69.780 75.850 69.805 ;
        RECT 82.210 69.780 82.560 69.805 ;
        RECT 88.920 69.780 89.270 69.805 ;
        RECT 95.630 69.780 95.980 69.805 ;
        RECT 102.340 69.780 102.690 69.805 ;
        RECT 105.345 69.790 105.675 69.805 ;
        RECT 37.560 69.355 37.910 69.380 ;
        RECT 44.270 69.355 44.620 69.380 ;
        RECT 37.560 69.055 44.620 69.355 ;
        RECT 37.560 69.030 37.910 69.055 ;
        RECT 44.270 69.030 44.620 69.055 ;
        RECT 50.980 69.355 51.330 69.380 ;
        RECT 57.690 69.355 58.040 69.380 ;
        RECT 50.980 69.055 58.040 69.355 ;
        RECT 50.980 69.030 51.330 69.055 ;
        RECT 57.690 69.030 58.040 69.055 ;
        RECT 64.400 69.355 64.750 69.380 ;
        RECT 71.110 69.355 71.460 69.380 ;
        RECT 64.400 69.055 71.460 69.355 ;
        RECT 64.400 69.030 64.750 69.055 ;
        RECT 71.110 69.030 71.460 69.055 ;
        RECT 77.820 69.355 78.170 69.380 ;
        RECT 84.530 69.355 84.880 69.380 ;
        RECT 77.820 69.055 84.880 69.355 ;
        RECT 77.820 69.030 78.170 69.055 ;
        RECT 84.530 69.030 84.880 69.055 ;
        RECT 91.240 69.355 91.590 69.380 ;
        RECT 97.950 69.355 98.300 69.380 ;
        RECT 91.240 69.055 98.300 69.355 ;
        RECT 91.240 69.030 91.590 69.055 ;
        RECT 97.950 69.030 98.300 69.055 ;
        RECT 33.305 68.605 33.635 68.620 ;
        RECT 36.290 68.605 36.640 68.630 ;
        RECT 43.000 68.605 43.350 68.630 ;
        RECT 49.710 68.605 50.060 68.630 ;
        RECT 56.420 68.605 56.770 68.630 ;
        RECT 63.130 68.605 63.480 68.630 ;
        RECT 69.840 68.605 70.190 68.630 ;
        RECT 76.550 68.605 76.900 68.630 ;
        RECT 83.260 68.605 83.610 68.630 ;
        RECT 89.970 68.605 90.320 68.630 ;
        RECT 96.680 68.605 97.030 68.630 ;
        RECT 106.845 68.605 107.175 68.620 ;
        RECT 33.305 68.305 107.175 68.605 ;
        RECT 33.305 68.290 33.635 68.305 ;
        RECT 36.290 68.280 36.640 68.305 ;
        RECT 43.000 68.280 43.350 68.305 ;
        RECT 49.710 68.280 50.060 68.305 ;
        RECT 56.420 68.280 56.770 68.305 ;
        RECT 63.130 68.280 63.480 68.305 ;
        RECT 69.840 68.280 70.190 68.305 ;
        RECT 76.550 68.280 76.900 68.305 ;
        RECT 83.260 68.280 83.610 68.305 ;
        RECT 89.970 68.280 90.320 68.305 ;
        RECT 96.680 68.280 97.030 68.305 ;
        RECT 106.845 68.290 107.175 68.305 ;
        RECT 37.980 67.855 38.330 67.880 ;
        RECT 44.690 67.855 45.040 67.880 ;
        RECT 37.980 67.555 45.040 67.855 ;
        RECT 37.980 67.530 38.330 67.555 ;
        RECT 44.690 67.530 45.040 67.555 ;
        RECT 51.400 67.855 51.750 67.880 ;
        RECT 58.110 67.855 58.460 67.880 ;
        RECT 51.400 67.555 58.460 67.855 ;
        RECT 51.400 67.530 51.750 67.555 ;
        RECT 58.110 67.530 58.460 67.555 ;
        RECT 64.820 67.855 65.170 67.880 ;
        RECT 71.530 67.855 71.880 67.880 ;
        RECT 64.820 67.555 71.880 67.855 ;
        RECT 64.820 67.530 65.170 67.555 ;
        RECT 71.530 67.530 71.880 67.555 ;
        RECT 78.240 67.855 78.590 67.880 ;
        RECT 84.950 67.855 85.300 67.880 ;
        RECT 78.240 67.555 85.300 67.855 ;
        RECT 78.240 67.530 78.590 67.555 ;
        RECT 84.950 67.530 85.300 67.555 ;
        RECT 91.660 67.855 92.010 67.880 ;
        RECT 98.370 67.855 98.720 67.880 ;
        RECT 91.660 67.555 98.720 67.855 ;
        RECT 91.660 67.530 92.010 67.555 ;
        RECT 98.370 67.530 98.720 67.555 ;
        RECT 34.805 67.105 35.135 67.120 ;
        RECT 41.950 67.105 42.300 67.130 ;
        RECT 48.660 67.105 49.010 67.130 ;
        RECT 55.370 67.105 55.720 67.130 ;
        RECT 62.080 67.105 62.430 67.130 ;
        RECT 68.790 67.105 69.140 67.130 ;
        RECT 75.500 67.105 75.850 67.130 ;
        RECT 82.210 67.105 82.560 67.130 ;
        RECT 88.920 67.105 89.270 67.130 ;
        RECT 95.630 67.105 95.980 67.130 ;
        RECT 102.340 67.105 102.690 67.130 ;
        RECT 105.345 67.105 105.675 67.120 ;
        RECT 34.805 66.805 105.675 67.105 ;
        RECT 34.805 66.790 35.135 66.805 ;
        RECT 41.950 66.780 42.300 66.805 ;
        RECT 48.660 66.780 49.010 66.805 ;
        RECT 55.370 66.780 55.720 66.805 ;
        RECT 62.080 66.780 62.430 66.805 ;
        RECT 68.790 66.780 69.140 66.805 ;
        RECT 75.500 66.780 75.850 66.805 ;
        RECT 82.210 66.780 82.560 66.805 ;
        RECT 88.920 66.780 89.270 66.805 ;
        RECT 95.630 66.780 95.980 66.805 ;
        RECT 102.340 66.780 102.690 66.805 ;
        RECT 105.345 66.790 105.675 66.805 ;
        RECT 37.140 66.355 37.490 66.380 ;
        RECT 43.850 66.355 44.200 66.380 ;
        RECT 37.140 66.055 44.200 66.355 ;
        RECT 37.140 66.030 37.490 66.055 ;
        RECT 43.850 66.030 44.200 66.055 ;
        RECT 50.560 66.355 50.910 66.380 ;
        RECT 57.270 66.355 57.620 66.380 ;
        RECT 50.560 66.055 57.620 66.355 ;
        RECT 50.560 66.030 50.910 66.055 ;
        RECT 57.270 66.030 57.620 66.055 ;
        RECT 63.980 66.355 64.330 66.380 ;
        RECT 70.690 66.355 71.040 66.380 ;
        RECT 63.980 66.055 71.040 66.355 ;
        RECT 63.980 66.030 64.330 66.055 ;
        RECT 70.690 66.030 71.040 66.055 ;
        RECT 77.400 66.355 77.750 66.380 ;
        RECT 84.110 66.355 84.460 66.380 ;
        RECT 77.400 66.055 84.460 66.355 ;
        RECT 77.400 66.030 77.750 66.055 ;
        RECT 84.110 66.030 84.460 66.055 ;
        RECT 90.820 66.355 91.170 66.380 ;
        RECT 97.530 66.355 97.880 66.380 ;
        RECT 90.820 66.055 97.880 66.355 ;
        RECT 90.820 66.030 91.170 66.055 ;
        RECT 97.530 66.030 97.880 66.055 ;
        RECT 33.305 65.605 33.635 65.620 ;
        RECT 36.290 65.605 36.640 65.630 ;
        RECT 43.000 65.605 43.350 65.630 ;
        RECT 49.710 65.605 50.060 65.630 ;
        RECT 56.420 65.605 56.770 65.630 ;
        RECT 63.130 65.605 63.480 65.630 ;
        RECT 69.840 65.605 70.190 65.630 ;
        RECT 76.550 65.605 76.900 65.630 ;
        RECT 83.260 65.605 83.610 65.630 ;
        RECT 89.970 65.605 90.320 65.630 ;
        RECT 96.680 65.605 97.030 65.630 ;
        RECT 101.500 65.605 101.830 65.620 ;
        RECT 106.845 65.605 107.175 65.620 ;
        RECT 33.305 65.305 107.175 65.605 ;
        RECT 33.305 65.290 33.635 65.305 ;
        RECT 36.290 65.280 36.640 65.305 ;
        RECT 43.000 65.280 43.350 65.305 ;
        RECT 49.710 65.280 50.060 65.305 ;
        RECT 56.420 65.280 56.770 65.305 ;
        RECT 63.130 65.280 63.480 65.305 ;
        RECT 69.840 65.280 70.190 65.305 ;
        RECT 76.550 65.280 76.900 65.305 ;
        RECT 83.260 65.280 83.610 65.305 ;
        RECT 89.970 65.280 90.320 65.305 ;
        RECT 96.680 65.280 97.030 65.305 ;
        RECT 101.500 65.290 101.830 65.305 ;
        RECT 106.845 65.290 107.175 65.305 ;
        RECT 38.500 63.735 39.500 63.765 ;
        RECT 71.500 63.735 72.500 63.765 ;
        RECT 104.500 63.735 105.500 63.765 ;
        RECT 30.325 62.735 108.305 63.735 ;
        RECT 38.500 62.715 39.500 62.735 ;
        RECT 71.500 62.715 72.500 62.735 ;
        RECT 104.500 62.715 105.500 62.735 ;
        RECT 35.500 61.735 36.500 61.765 ;
        RECT 68.500 61.735 69.500 61.765 ;
        RECT 101.500 61.735 102.500 61.765 ;
        RECT 30.325 60.735 108.305 61.735 ;
        RECT 35.500 60.715 36.500 60.735 ;
        RECT 68.500 60.715 69.500 60.735 ;
        RECT 101.500 60.715 102.500 60.735 ;
        RECT 110.325 59.925 110.625 184.700 ;
        RECT 110.955 60.335 111.255 185.700 ;
        RECT 110.940 60.005 111.270 60.335 ;
        RECT 32.500 59.735 33.500 59.765 ;
        RECT 65.500 59.735 66.500 59.765 ;
        RECT 98.500 59.735 99.500 59.765 ;
        RECT 30.325 58.735 108.305 59.735 ;
        RECT 110.310 59.595 110.640 59.925 ;
        RECT 111.585 59.105 111.885 186.700 ;
        RECT 112.215 186.700 112.980 187.000 ;
        RECT 112.215 164.705 112.515 186.700 ;
        RECT 114.180 186.000 114.480 189.015 ;
        RECT 112.845 185.700 114.480 186.000 ;
        RECT 112.845 165.525 113.145 185.700 ;
        RECT 115.680 185.000 115.980 189.015 ;
        RECT 113.475 184.700 115.980 185.000 ;
        RECT 113.475 165.935 113.775 184.700 ;
        RECT 117.180 184.020 117.480 189.015 ;
        RECT 114.105 183.720 117.480 184.020 ;
        RECT 113.460 165.605 113.790 165.935 ;
        RECT 112.830 165.195 113.160 165.525 ;
        RECT 112.200 164.375 112.530 164.705 ;
        RECT 112.215 59.515 112.515 164.375 ;
        RECT 112.845 60.735 113.145 165.195 ;
        RECT 114.105 164.295 114.405 183.720 ;
        RECT 117.180 183.700 117.480 183.720 ;
        RECT 118.680 183.000 118.980 189.015 ;
        RECT 114.735 182.700 118.980 183.000 ;
        RECT 114.735 165.115 115.035 182.700 ;
        RECT 114.720 164.785 115.050 165.115 ;
        RECT 114.090 163.965 114.420 164.295 ;
        RECT 115.060 129.625 137.070 130.525 ;
        RECT 112.200 59.185 112.530 59.515 ;
        RECT 111.570 58.775 111.900 59.105 ;
        RECT 32.500 58.715 33.500 58.735 ;
        RECT 65.500 58.715 66.500 58.735 ;
        RECT 98.500 58.715 99.500 58.735 ;
        RECT 136.170 0.995 137.070 129.625 ;
        RECT 136.145 0.105 137.095 0.995 ;
        RECT 136.170 0.100 137.070 0.105 ;
      LAYER met4 ;
        RECT 15.015 224.760 15.030 225.075 ;
        RECT 15.330 224.760 15.345 225.075 ;
        RECT 15.015 224.745 15.345 224.760 ;
        RECT 17.775 224.760 17.790 225.075 ;
        RECT 18.090 224.760 18.105 225.075 ;
        RECT 17.775 224.745 18.105 224.760 ;
        RECT 20.535 224.760 20.550 225.075 ;
        RECT 20.850 224.760 20.865 225.075 ;
        RECT 20.535 224.745 20.865 224.760 ;
        RECT 23.295 224.760 23.310 225.075 ;
        RECT 23.610 224.760 23.625 225.075 ;
        RECT 23.295 224.745 23.625 224.760 ;
        RECT 26.055 224.760 26.070 225.075 ;
        RECT 26.370 224.760 26.385 225.075 ;
        RECT 26.055 224.745 26.385 224.760 ;
        RECT 28.815 224.760 28.830 225.075 ;
        RECT 29.130 224.760 29.145 225.075 ;
        RECT 28.815 224.745 29.145 224.760 ;
        RECT 31.575 224.760 31.590 225.075 ;
        RECT 31.890 224.760 31.905 225.075 ;
        RECT 31.575 224.745 31.905 224.760 ;
        RECT 34.335 224.760 34.350 225.075 ;
        RECT 34.650 224.760 34.665 225.075 ;
        RECT 34.335 224.745 34.665 224.760 ;
        RECT 37.095 224.760 37.110 225.075 ;
        RECT 37.410 224.760 37.425 225.075 ;
        RECT 37.095 224.745 37.425 224.760 ;
        RECT 39.855 224.760 39.870 225.075 ;
        RECT 40.170 224.760 40.185 225.075 ;
        RECT 39.855 224.745 40.185 224.760 ;
        RECT 42.615 224.760 42.630 225.075 ;
        RECT 42.930 224.760 42.945 225.075 ;
        RECT 42.615 224.745 42.945 224.760 ;
        RECT 45.375 224.760 45.390 225.075 ;
        RECT 45.690 224.760 45.705 225.075 ;
        RECT 45.375 224.745 45.705 224.760 ;
        RECT 48.135 224.760 48.150 225.075 ;
        RECT 48.450 224.760 48.465 225.075 ;
        RECT 48.135 224.745 48.465 224.760 ;
        RECT 50.895 224.760 50.910 225.075 ;
        RECT 51.210 224.760 51.225 225.075 ;
        RECT 50.895 224.745 51.225 224.760 ;
        RECT 53.655 224.760 53.670 225.075 ;
        RECT 53.970 224.760 53.985 225.075 ;
        RECT 53.655 224.745 53.985 224.760 ;
        RECT 56.415 224.760 56.430 225.075 ;
        RECT 56.730 224.760 56.745 225.075 ;
        RECT 56.415 224.745 56.745 224.760 ;
        RECT 59.175 224.760 59.190 225.075 ;
        RECT 59.490 224.760 59.505 225.075 ;
        RECT 59.175 224.745 59.505 224.760 ;
        RECT 61.935 224.760 61.950 225.075 ;
        RECT 62.250 224.760 62.265 225.075 ;
        RECT 61.935 224.745 62.265 224.760 ;
        RECT 64.695 224.760 64.710 225.075 ;
        RECT 65.010 224.760 65.025 225.075 ;
        RECT 64.695 224.745 65.025 224.760 ;
        RECT 67.455 224.760 67.470 225.075 ;
        RECT 67.770 224.760 67.785 225.075 ;
        RECT 67.455 224.745 67.785 224.760 ;
        RECT 70.215 224.760 70.230 225.075 ;
        RECT 70.530 224.760 70.545 225.075 ;
        RECT 70.215 224.745 70.545 224.760 ;
        RECT 72.975 224.760 72.990 225.075 ;
        RECT 73.290 224.760 73.305 225.075 ;
        RECT 72.975 224.745 73.305 224.760 ;
        RECT 75.735 224.760 75.750 225.075 ;
        RECT 76.050 224.760 76.065 225.075 ;
        RECT 75.735 224.745 76.065 224.760 ;
        RECT 78.495 224.760 78.510 225.075 ;
        RECT 78.810 224.760 78.825 225.075 ;
        RECT 78.495 224.745 78.825 224.760 ;
        RECT 103.335 224.760 103.350 225.075 ;
        RECT 103.650 224.760 103.665 225.075 ;
        RECT 103.335 224.745 103.665 224.760 ;
        RECT 106.095 224.760 106.110 225.075 ;
        RECT 106.410 224.760 106.425 225.075 ;
        RECT 106.095 224.745 106.425 224.760 ;
        RECT 108.855 224.760 108.870 225.075 ;
        RECT 109.170 224.760 109.185 225.075 ;
        RECT 108.855 224.745 109.185 224.760 ;
        RECT 111.615 224.760 111.630 225.075 ;
        RECT 111.930 224.760 111.945 225.075 ;
        RECT 111.615 224.745 111.945 224.760 ;
        RECT 114.375 224.760 114.390 225.075 ;
        RECT 114.690 224.760 114.705 225.075 ;
        RECT 114.375 224.745 114.705 224.760 ;
        RECT 117.135 224.760 117.150 225.075 ;
        RECT 117.450 224.760 117.465 225.075 ;
        RECT 117.135 224.745 117.465 224.760 ;
        RECT 119.895 224.760 119.910 225.085 ;
        RECT 120.210 224.760 120.225 225.085 ;
        RECT 119.895 224.755 120.225 224.760 ;
        RECT 122.655 224.760 122.670 225.075 ;
        RECT 122.970 224.760 122.985 225.075 ;
        RECT 122.655 224.745 122.985 224.760 ;
  END
END tt_um_htfab_dg_dac
END LIBRARY

